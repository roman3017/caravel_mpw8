VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO user_proj_example
  CLASS BLOCK ;
  FOREIGN user_proj_example ;
  ORIGIN 0.000 0.000 ;
  SIZE 900.000 BY 600.000 ;
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 7.910 596.000 8.190 600.000 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 242.510 596.000 242.790 600.000 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 265.970 596.000 266.250 600.000 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 289.430 596.000 289.710 600.000 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 312.890 596.000 313.170 600.000 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 336.350 596.000 336.630 600.000 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 359.810 596.000 360.090 600.000 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 383.270 596.000 383.550 600.000 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 406.730 596.000 407.010 600.000 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 430.190 596.000 430.470 600.000 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 453.650 596.000 453.930 600.000 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 31.370 596.000 31.650 600.000 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 477.110 596.000 477.390 600.000 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 500.570 596.000 500.850 600.000 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 524.030 596.000 524.310 600.000 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 547.490 596.000 547.770 600.000 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 570.950 596.000 571.230 600.000 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 594.410 596.000 594.690 600.000 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 617.870 596.000 618.150 600.000 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 641.330 596.000 641.610 600.000 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 664.790 596.000 665.070 600.000 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 688.250 596.000 688.530 600.000 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.830 596.000 55.110 600.000 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 711.710 596.000 711.990 600.000 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 735.170 596.000 735.450 600.000 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 758.630 596.000 758.910 600.000 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 782.090 596.000 782.370 600.000 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 805.550 596.000 805.830 600.000 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 829.010 596.000 829.290 600.000 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 852.470 596.000 852.750 600.000 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 875.930 596.000 876.210 600.000 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 78.290 596.000 78.570 600.000 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 101.750 596.000 102.030 600.000 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 125.210 596.000 125.490 600.000 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 148.670 596.000 148.950 600.000 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 172.130 596.000 172.410 600.000 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 195.590 596.000 195.870 600.000 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 219.050 596.000 219.330 600.000 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 15.730 596.000 16.010 600.000 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 250.330 596.000 250.610 600.000 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 273.790 596.000 274.070 600.000 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 297.250 596.000 297.530 600.000 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 320.710 596.000 320.990 600.000 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 344.170 596.000 344.450 600.000 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 367.630 596.000 367.910 600.000 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 391.090 596.000 391.370 600.000 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 414.550 596.000 414.830 600.000 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 438.010 596.000 438.290 600.000 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 461.470 596.000 461.750 600.000 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.190 596.000 39.470 600.000 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 484.930 596.000 485.210 600.000 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 508.390 596.000 508.670 600.000 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 531.850 596.000 532.130 600.000 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 555.310 596.000 555.590 600.000 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 578.770 596.000 579.050 600.000 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 602.230 596.000 602.510 600.000 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 625.690 596.000 625.970 600.000 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 649.150 596.000 649.430 600.000 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 672.610 596.000 672.890 600.000 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 696.070 596.000 696.350 600.000 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.650 596.000 62.930 600.000 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 719.530 596.000 719.810 600.000 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 742.990 596.000 743.270 600.000 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 766.450 596.000 766.730 600.000 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 789.910 596.000 790.190 600.000 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 813.370 596.000 813.650 600.000 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 836.830 596.000 837.110 600.000 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 860.290 596.000 860.570 600.000 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 883.750 596.000 884.030 600.000 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 86.110 596.000 86.390 600.000 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.570 596.000 109.850 600.000 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 133.030 596.000 133.310 600.000 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 156.490 596.000 156.770 600.000 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 179.950 596.000 180.230 600.000 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 203.410 596.000 203.690 600.000 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 226.870 596.000 227.150 600.000 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 23.550 596.000 23.830 600.000 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 258.150 596.000 258.430 600.000 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 281.610 596.000 281.890 600.000 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 305.070 596.000 305.350 600.000 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 328.530 596.000 328.810 600.000 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 351.990 596.000 352.270 600.000 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 375.450 596.000 375.730 600.000 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 398.910 596.000 399.190 600.000 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 422.370 596.000 422.650 600.000 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 445.830 596.000 446.110 600.000 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 469.290 596.000 469.570 600.000 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.010 596.000 47.290 600.000 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 492.750 596.000 493.030 600.000 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 516.210 596.000 516.490 600.000 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 539.670 596.000 539.950 600.000 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 563.130 596.000 563.410 600.000 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 586.590 596.000 586.870 600.000 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 610.050 596.000 610.330 600.000 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 633.510 596.000 633.790 600.000 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 656.970 596.000 657.250 600.000 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 680.430 596.000 680.710 600.000 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 703.890 596.000 704.170 600.000 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.470 596.000 70.750 600.000 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 727.350 596.000 727.630 600.000 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 750.810 596.000 751.090 600.000 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 774.270 596.000 774.550 600.000 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 797.730 596.000 798.010 600.000 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 821.190 596.000 821.470 600.000 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 844.650 596.000 844.930 600.000 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 868.110 596.000 868.390 600.000 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 891.570 596.000 891.850 600.000 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.930 596.000 94.210 600.000 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 117.390 596.000 117.670 600.000 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 140.850 596.000 141.130 600.000 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 164.310 596.000 164.590 600.000 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 187.770 596.000 188.050 600.000 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 211.230 596.000 211.510 600.000 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 234.690 596.000 234.970 600.000 ;
    END
  END io_out[9]
  PIN irq[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 787.150 0.000 787.430 4.000 ;
    END
  END irq[0]
  PIN irq[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 788.530 0.000 788.810 4.000 ;
    END
  END irq[1]
  PIN irq[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 789.910 0.000 790.190 4.000 ;
    END
  END irq[2]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 255.850 0.000 256.130 4.000 ;
    END
  END la_data_in[0]
  PIN la_data_in[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 669.850 0.000 670.130 4.000 ;
    END
  END la_data_in[100]
  PIN la_data_in[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 673.990 0.000 674.270 4.000 ;
    END
  END la_data_in[101]
  PIN la_data_in[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 678.130 0.000 678.410 4.000 ;
    END
  END la_data_in[102]
  PIN la_data_in[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 682.270 0.000 682.550 4.000 ;
    END
  END la_data_in[103]
  PIN la_data_in[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 686.410 0.000 686.690 4.000 ;
    END
  END la_data_in[104]
  PIN la_data_in[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 690.550 0.000 690.830 4.000 ;
    END
  END la_data_in[105]
  PIN la_data_in[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 694.690 0.000 694.970 4.000 ;
    END
  END la_data_in[106]
  PIN la_data_in[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 698.830 0.000 699.110 4.000 ;
    END
  END la_data_in[107]
  PIN la_data_in[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 702.970 0.000 703.250 4.000 ;
    END
  END la_data_in[108]
  PIN la_data_in[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 707.110 0.000 707.390 4.000 ;
    END
  END la_data_in[109]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 297.250 0.000 297.530 4.000 ;
    END
  END la_data_in[10]
  PIN la_data_in[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 711.250 0.000 711.530 4.000 ;
    END
  END la_data_in[110]
  PIN la_data_in[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 715.390 0.000 715.670 4.000 ;
    END
  END la_data_in[111]
  PIN la_data_in[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 719.530 0.000 719.810 4.000 ;
    END
  END la_data_in[112]
  PIN la_data_in[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 723.670 0.000 723.950 4.000 ;
    END
  END la_data_in[113]
  PIN la_data_in[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 727.810 0.000 728.090 4.000 ;
    END
  END la_data_in[114]
  PIN la_data_in[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 731.950 0.000 732.230 4.000 ;
    END
  END la_data_in[115]
  PIN la_data_in[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 736.090 0.000 736.370 4.000 ;
    END
  END la_data_in[116]
  PIN la_data_in[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 740.230 0.000 740.510 4.000 ;
    END
  END la_data_in[117]
  PIN la_data_in[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 744.370 0.000 744.650 4.000 ;
    END
  END la_data_in[118]
  PIN la_data_in[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 748.510 0.000 748.790 4.000 ;
    END
  END la_data_in[119]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 301.390 0.000 301.670 4.000 ;
    END
  END la_data_in[11]
  PIN la_data_in[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 752.650 0.000 752.930 4.000 ;
    END
  END la_data_in[120]
  PIN la_data_in[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 756.790 0.000 757.070 4.000 ;
    END
  END la_data_in[121]
  PIN la_data_in[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 760.930 0.000 761.210 4.000 ;
    END
  END la_data_in[122]
  PIN la_data_in[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 765.070 0.000 765.350 4.000 ;
    END
  END la_data_in[123]
  PIN la_data_in[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 769.210 0.000 769.490 4.000 ;
    END
  END la_data_in[124]
  PIN la_data_in[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 773.350 0.000 773.630 4.000 ;
    END
  END la_data_in[125]
  PIN la_data_in[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 777.490 0.000 777.770 4.000 ;
    END
  END la_data_in[126]
  PIN la_data_in[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 781.630 0.000 781.910 4.000 ;
    END
  END la_data_in[127]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 305.530 0.000 305.810 4.000 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 309.670 0.000 309.950 4.000 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 313.810 0.000 314.090 4.000 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 317.950 0.000 318.230 4.000 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 322.090 0.000 322.370 4.000 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 326.230 0.000 326.510 4.000 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 330.370 0.000 330.650 4.000 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 334.510 0.000 334.790 4.000 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 259.990 0.000 260.270 4.000 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 338.650 0.000 338.930 4.000 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 342.790 0.000 343.070 4.000 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 346.930 0.000 347.210 4.000 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 351.070 0.000 351.350 4.000 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 355.210 0.000 355.490 4.000 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 359.350 0.000 359.630 4.000 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 363.490 0.000 363.770 4.000 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 367.630 0.000 367.910 4.000 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 371.770 0.000 372.050 4.000 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 375.910 0.000 376.190 4.000 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 264.130 0.000 264.410 4.000 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 380.050 0.000 380.330 4.000 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 384.190 0.000 384.470 4.000 ;
    END
  END la_data_in[31]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 388.330 0.000 388.610 4.000 ;
    END
  END la_data_in[32]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 392.470 0.000 392.750 4.000 ;
    END
  END la_data_in[33]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 396.610 0.000 396.890 4.000 ;
    END
  END la_data_in[34]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 400.750 0.000 401.030 4.000 ;
    END
  END la_data_in[35]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 404.890 0.000 405.170 4.000 ;
    END
  END la_data_in[36]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 409.030 0.000 409.310 4.000 ;
    END
  END la_data_in[37]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 413.170 0.000 413.450 4.000 ;
    END
  END la_data_in[38]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 417.310 0.000 417.590 4.000 ;
    END
  END la_data_in[39]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 268.270 0.000 268.550 4.000 ;
    END
  END la_data_in[3]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 421.450 0.000 421.730 4.000 ;
    END
  END la_data_in[40]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 425.590 0.000 425.870 4.000 ;
    END
  END la_data_in[41]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 429.730 0.000 430.010 4.000 ;
    END
  END la_data_in[42]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 433.870 0.000 434.150 4.000 ;
    END
  END la_data_in[43]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 438.010 0.000 438.290 4.000 ;
    END
  END la_data_in[44]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 442.150 0.000 442.430 4.000 ;
    END
  END la_data_in[45]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 446.290 0.000 446.570 4.000 ;
    END
  END la_data_in[46]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 450.430 0.000 450.710 4.000 ;
    END
  END la_data_in[47]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 454.570 0.000 454.850 4.000 ;
    END
  END la_data_in[48]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 458.710 0.000 458.990 4.000 ;
    END
  END la_data_in[49]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 272.410 0.000 272.690 4.000 ;
    END
  END la_data_in[4]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 462.850 0.000 463.130 4.000 ;
    END
  END la_data_in[50]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 466.990 0.000 467.270 4.000 ;
    END
  END la_data_in[51]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 471.130 0.000 471.410 4.000 ;
    END
  END la_data_in[52]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 475.270 0.000 475.550 4.000 ;
    END
  END la_data_in[53]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 479.410 0.000 479.690 4.000 ;
    END
  END la_data_in[54]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 483.550 0.000 483.830 4.000 ;
    END
  END la_data_in[55]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 487.690 0.000 487.970 4.000 ;
    END
  END la_data_in[56]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 491.830 0.000 492.110 4.000 ;
    END
  END la_data_in[57]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 495.970 0.000 496.250 4.000 ;
    END
  END la_data_in[58]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 500.110 0.000 500.390 4.000 ;
    END
  END la_data_in[59]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 276.550 0.000 276.830 4.000 ;
    END
  END la_data_in[5]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 504.250 0.000 504.530 4.000 ;
    END
  END la_data_in[60]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 508.390 0.000 508.670 4.000 ;
    END
  END la_data_in[61]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 512.530 0.000 512.810 4.000 ;
    END
  END la_data_in[62]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 516.670 0.000 516.950 4.000 ;
    END
  END la_data_in[63]
  PIN la_data_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 520.810 0.000 521.090 4.000 ;
    END
  END la_data_in[64]
  PIN la_data_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 524.950 0.000 525.230 4.000 ;
    END
  END la_data_in[65]
  PIN la_data_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 529.090 0.000 529.370 4.000 ;
    END
  END la_data_in[66]
  PIN la_data_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 533.230 0.000 533.510 4.000 ;
    END
  END la_data_in[67]
  PIN la_data_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 537.370 0.000 537.650 4.000 ;
    END
  END la_data_in[68]
  PIN la_data_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 541.510 0.000 541.790 4.000 ;
    END
  END la_data_in[69]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 280.690 0.000 280.970 4.000 ;
    END
  END la_data_in[6]
  PIN la_data_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 545.650 0.000 545.930 4.000 ;
    END
  END la_data_in[70]
  PIN la_data_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 549.790 0.000 550.070 4.000 ;
    END
  END la_data_in[71]
  PIN la_data_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 553.930 0.000 554.210 4.000 ;
    END
  END la_data_in[72]
  PIN la_data_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 558.070 0.000 558.350 4.000 ;
    END
  END la_data_in[73]
  PIN la_data_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 562.210 0.000 562.490 4.000 ;
    END
  END la_data_in[74]
  PIN la_data_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 566.350 0.000 566.630 4.000 ;
    END
  END la_data_in[75]
  PIN la_data_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 570.490 0.000 570.770 4.000 ;
    END
  END la_data_in[76]
  PIN la_data_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 574.630 0.000 574.910 4.000 ;
    END
  END la_data_in[77]
  PIN la_data_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 578.770 0.000 579.050 4.000 ;
    END
  END la_data_in[78]
  PIN la_data_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 582.910 0.000 583.190 4.000 ;
    END
  END la_data_in[79]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 284.830 0.000 285.110 4.000 ;
    END
  END la_data_in[7]
  PIN la_data_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 587.050 0.000 587.330 4.000 ;
    END
  END la_data_in[80]
  PIN la_data_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 591.190 0.000 591.470 4.000 ;
    END
  END la_data_in[81]
  PIN la_data_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 595.330 0.000 595.610 4.000 ;
    END
  END la_data_in[82]
  PIN la_data_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 599.470 0.000 599.750 4.000 ;
    END
  END la_data_in[83]
  PIN la_data_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 603.610 0.000 603.890 4.000 ;
    END
  END la_data_in[84]
  PIN la_data_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 607.750 0.000 608.030 4.000 ;
    END
  END la_data_in[85]
  PIN la_data_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 611.890 0.000 612.170 4.000 ;
    END
  END la_data_in[86]
  PIN la_data_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 616.030 0.000 616.310 4.000 ;
    END
  END la_data_in[87]
  PIN la_data_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 620.170 0.000 620.450 4.000 ;
    END
  END la_data_in[88]
  PIN la_data_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 624.310 0.000 624.590 4.000 ;
    END
  END la_data_in[89]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 288.970 0.000 289.250 4.000 ;
    END
  END la_data_in[8]
  PIN la_data_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 628.450 0.000 628.730 4.000 ;
    END
  END la_data_in[90]
  PIN la_data_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 632.590 0.000 632.870 4.000 ;
    END
  END la_data_in[91]
  PIN la_data_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 636.730 0.000 637.010 4.000 ;
    END
  END la_data_in[92]
  PIN la_data_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 640.870 0.000 641.150 4.000 ;
    END
  END la_data_in[93]
  PIN la_data_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 645.010 0.000 645.290 4.000 ;
    END
  END la_data_in[94]
  PIN la_data_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 649.150 0.000 649.430 4.000 ;
    END
  END la_data_in[95]
  PIN la_data_in[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 653.290 0.000 653.570 4.000 ;
    END
  END la_data_in[96]
  PIN la_data_in[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 657.430 0.000 657.710 4.000 ;
    END
  END la_data_in[97]
  PIN la_data_in[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 661.570 0.000 661.850 4.000 ;
    END
  END la_data_in[98]
  PIN la_data_in[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 665.710 0.000 665.990 4.000 ;
    END
  END la_data_in[99]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 293.110 0.000 293.390 4.000 ;
    END
  END la_data_in[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 257.230 0.000 257.510 4.000 ;
    END
  END la_data_out[0]
  PIN la_data_out[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 671.230 0.000 671.510 4.000 ;
    END
  END la_data_out[100]
  PIN la_data_out[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 675.370 0.000 675.650 4.000 ;
    END
  END la_data_out[101]
  PIN la_data_out[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 679.510 0.000 679.790 4.000 ;
    END
  END la_data_out[102]
  PIN la_data_out[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 683.650 0.000 683.930 4.000 ;
    END
  END la_data_out[103]
  PIN la_data_out[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 687.790 0.000 688.070 4.000 ;
    END
  END la_data_out[104]
  PIN la_data_out[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 691.930 0.000 692.210 4.000 ;
    END
  END la_data_out[105]
  PIN la_data_out[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 696.070 0.000 696.350 4.000 ;
    END
  END la_data_out[106]
  PIN la_data_out[107]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 700.210 0.000 700.490 4.000 ;
    END
  END la_data_out[107]
  PIN la_data_out[108]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 704.350 0.000 704.630 4.000 ;
    END
  END la_data_out[108]
  PIN la_data_out[109]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 708.490 0.000 708.770 4.000 ;
    END
  END la_data_out[109]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 298.630 0.000 298.910 4.000 ;
    END
  END la_data_out[10]
  PIN la_data_out[110]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 712.630 0.000 712.910 4.000 ;
    END
  END la_data_out[110]
  PIN la_data_out[111]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 716.770 0.000 717.050 4.000 ;
    END
  END la_data_out[111]
  PIN la_data_out[112]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 720.910 0.000 721.190 4.000 ;
    END
  END la_data_out[112]
  PIN la_data_out[113]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 725.050 0.000 725.330 4.000 ;
    END
  END la_data_out[113]
  PIN la_data_out[114]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 729.190 0.000 729.470 4.000 ;
    END
  END la_data_out[114]
  PIN la_data_out[115]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 733.330 0.000 733.610 4.000 ;
    END
  END la_data_out[115]
  PIN la_data_out[116]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 737.470 0.000 737.750 4.000 ;
    END
  END la_data_out[116]
  PIN la_data_out[117]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 741.610 0.000 741.890 4.000 ;
    END
  END la_data_out[117]
  PIN la_data_out[118]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 745.750 0.000 746.030 4.000 ;
    END
  END la_data_out[118]
  PIN la_data_out[119]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 749.890 0.000 750.170 4.000 ;
    END
  END la_data_out[119]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 302.770 0.000 303.050 4.000 ;
    END
  END la_data_out[11]
  PIN la_data_out[120]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 754.030 0.000 754.310 4.000 ;
    END
  END la_data_out[120]
  PIN la_data_out[121]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 758.170 0.000 758.450 4.000 ;
    END
  END la_data_out[121]
  PIN la_data_out[122]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 762.310 0.000 762.590 4.000 ;
    END
  END la_data_out[122]
  PIN la_data_out[123]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 766.450 0.000 766.730 4.000 ;
    END
  END la_data_out[123]
  PIN la_data_out[124]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 770.590 0.000 770.870 4.000 ;
    END
  END la_data_out[124]
  PIN la_data_out[125]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 774.730 0.000 775.010 4.000 ;
    END
  END la_data_out[125]
  PIN la_data_out[126]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 778.870 0.000 779.150 4.000 ;
    END
  END la_data_out[126]
  PIN la_data_out[127]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 783.010 0.000 783.290 4.000 ;
    END
  END la_data_out[127]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 306.910 0.000 307.190 4.000 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 311.050 0.000 311.330 4.000 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 315.190 0.000 315.470 4.000 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 319.330 0.000 319.610 4.000 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 323.470 0.000 323.750 4.000 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 327.610 0.000 327.890 4.000 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 331.750 0.000 332.030 4.000 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 335.890 0.000 336.170 4.000 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 261.370 0.000 261.650 4.000 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 340.030 0.000 340.310 4.000 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 344.170 0.000 344.450 4.000 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 348.310 0.000 348.590 4.000 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 352.450 0.000 352.730 4.000 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 356.590 0.000 356.870 4.000 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 360.730 0.000 361.010 4.000 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 364.870 0.000 365.150 4.000 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 369.010 0.000 369.290 4.000 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 373.150 0.000 373.430 4.000 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 377.290 0.000 377.570 4.000 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 265.510 0.000 265.790 4.000 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 381.430 0.000 381.710 4.000 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 385.570 0.000 385.850 4.000 ;
    END
  END la_data_out[31]
  PIN la_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 389.710 0.000 389.990 4.000 ;
    END
  END la_data_out[32]
  PIN la_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 393.850 0.000 394.130 4.000 ;
    END
  END la_data_out[33]
  PIN la_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 397.990 0.000 398.270 4.000 ;
    END
  END la_data_out[34]
  PIN la_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 402.130 0.000 402.410 4.000 ;
    END
  END la_data_out[35]
  PIN la_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 406.270 0.000 406.550 4.000 ;
    END
  END la_data_out[36]
  PIN la_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 410.410 0.000 410.690 4.000 ;
    END
  END la_data_out[37]
  PIN la_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 414.550 0.000 414.830 4.000 ;
    END
  END la_data_out[38]
  PIN la_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 418.690 0.000 418.970 4.000 ;
    END
  END la_data_out[39]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 269.650 0.000 269.930 4.000 ;
    END
  END la_data_out[3]
  PIN la_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 422.830 0.000 423.110 4.000 ;
    END
  END la_data_out[40]
  PIN la_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 426.970 0.000 427.250 4.000 ;
    END
  END la_data_out[41]
  PIN la_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 431.110 0.000 431.390 4.000 ;
    END
  END la_data_out[42]
  PIN la_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 435.250 0.000 435.530 4.000 ;
    END
  END la_data_out[43]
  PIN la_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 439.390 0.000 439.670 4.000 ;
    END
  END la_data_out[44]
  PIN la_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 443.530 0.000 443.810 4.000 ;
    END
  END la_data_out[45]
  PIN la_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 447.670 0.000 447.950 4.000 ;
    END
  END la_data_out[46]
  PIN la_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 451.810 0.000 452.090 4.000 ;
    END
  END la_data_out[47]
  PIN la_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 455.950 0.000 456.230 4.000 ;
    END
  END la_data_out[48]
  PIN la_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 460.090 0.000 460.370 4.000 ;
    END
  END la_data_out[49]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 273.790 0.000 274.070 4.000 ;
    END
  END la_data_out[4]
  PIN la_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 464.230 0.000 464.510 4.000 ;
    END
  END la_data_out[50]
  PIN la_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 468.370 0.000 468.650 4.000 ;
    END
  END la_data_out[51]
  PIN la_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 472.510 0.000 472.790 4.000 ;
    END
  END la_data_out[52]
  PIN la_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 476.650 0.000 476.930 4.000 ;
    END
  END la_data_out[53]
  PIN la_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 480.790 0.000 481.070 4.000 ;
    END
  END la_data_out[54]
  PIN la_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 484.930 0.000 485.210 4.000 ;
    END
  END la_data_out[55]
  PIN la_data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 489.070 0.000 489.350 4.000 ;
    END
  END la_data_out[56]
  PIN la_data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 493.210 0.000 493.490 4.000 ;
    END
  END la_data_out[57]
  PIN la_data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 497.350 0.000 497.630 4.000 ;
    END
  END la_data_out[58]
  PIN la_data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 501.490 0.000 501.770 4.000 ;
    END
  END la_data_out[59]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 277.930 0.000 278.210 4.000 ;
    END
  END la_data_out[5]
  PIN la_data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 505.630 0.000 505.910 4.000 ;
    END
  END la_data_out[60]
  PIN la_data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 509.770 0.000 510.050 4.000 ;
    END
  END la_data_out[61]
  PIN la_data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 513.910 0.000 514.190 4.000 ;
    END
  END la_data_out[62]
  PIN la_data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 518.050 0.000 518.330 4.000 ;
    END
  END la_data_out[63]
  PIN la_data_out[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 522.190 0.000 522.470 4.000 ;
    END
  END la_data_out[64]
  PIN la_data_out[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 526.330 0.000 526.610 4.000 ;
    END
  END la_data_out[65]
  PIN la_data_out[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 530.470 0.000 530.750 4.000 ;
    END
  END la_data_out[66]
  PIN la_data_out[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 534.610 0.000 534.890 4.000 ;
    END
  END la_data_out[67]
  PIN la_data_out[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 538.750 0.000 539.030 4.000 ;
    END
  END la_data_out[68]
  PIN la_data_out[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 542.890 0.000 543.170 4.000 ;
    END
  END la_data_out[69]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 282.070 0.000 282.350 4.000 ;
    END
  END la_data_out[6]
  PIN la_data_out[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 547.030 0.000 547.310 4.000 ;
    END
  END la_data_out[70]
  PIN la_data_out[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 551.170 0.000 551.450 4.000 ;
    END
  END la_data_out[71]
  PIN la_data_out[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 555.310 0.000 555.590 4.000 ;
    END
  END la_data_out[72]
  PIN la_data_out[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 559.450 0.000 559.730 4.000 ;
    END
  END la_data_out[73]
  PIN la_data_out[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 563.590 0.000 563.870 4.000 ;
    END
  END la_data_out[74]
  PIN la_data_out[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 567.730 0.000 568.010 4.000 ;
    END
  END la_data_out[75]
  PIN la_data_out[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 571.870 0.000 572.150 4.000 ;
    END
  END la_data_out[76]
  PIN la_data_out[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 576.010 0.000 576.290 4.000 ;
    END
  END la_data_out[77]
  PIN la_data_out[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 580.150 0.000 580.430 4.000 ;
    END
  END la_data_out[78]
  PIN la_data_out[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 584.290 0.000 584.570 4.000 ;
    END
  END la_data_out[79]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 286.210 0.000 286.490 4.000 ;
    END
  END la_data_out[7]
  PIN la_data_out[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 588.430 0.000 588.710 4.000 ;
    END
  END la_data_out[80]
  PIN la_data_out[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 592.570 0.000 592.850 4.000 ;
    END
  END la_data_out[81]
  PIN la_data_out[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 596.710 0.000 596.990 4.000 ;
    END
  END la_data_out[82]
  PIN la_data_out[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 600.850 0.000 601.130 4.000 ;
    END
  END la_data_out[83]
  PIN la_data_out[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 604.990 0.000 605.270 4.000 ;
    END
  END la_data_out[84]
  PIN la_data_out[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 609.130 0.000 609.410 4.000 ;
    END
  END la_data_out[85]
  PIN la_data_out[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 613.270 0.000 613.550 4.000 ;
    END
  END la_data_out[86]
  PIN la_data_out[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 617.410 0.000 617.690 4.000 ;
    END
  END la_data_out[87]
  PIN la_data_out[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 621.550 0.000 621.830 4.000 ;
    END
  END la_data_out[88]
  PIN la_data_out[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 625.690 0.000 625.970 4.000 ;
    END
  END la_data_out[89]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 290.350 0.000 290.630 4.000 ;
    END
  END la_data_out[8]
  PIN la_data_out[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 629.830 0.000 630.110 4.000 ;
    END
  END la_data_out[90]
  PIN la_data_out[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 633.970 0.000 634.250 4.000 ;
    END
  END la_data_out[91]
  PIN la_data_out[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 638.110 0.000 638.390 4.000 ;
    END
  END la_data_out[92]
  PIN la_data_out[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 642.250 0.000 642.530 4.000 ;
    END
  END la_data_out[93]
  PIN la_data_out[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 646.390 0.000 646.670 4.000 ;
    END
  END la_data_out[94]
  PIN la_data_out[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 650.530 0.000 650.810 4.000 ;
    END
  END la_data_out[95]
  PIN la_data_out[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 654.670 0.000 654.950 4.000 ;
    END
  END la_data_out[96]
  PIN la_data_out[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 658.810 0.000 659.090 4.000 ;
    END
  END la_data_out[97]
  PIN la_data_out[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 662.950 0.000 663.230 4.000 ;
    END
  END la_data_out[98]
  PIN la_data_out[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 667.090 0.000 667.370 4.000 ;
    END
  END la_data_out[99]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 294.490 0.000 294.770 4.000 ;
    END
  END la_data_out[9]
  PIN la_oenb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 258.610 0.000 258.890 4.000 ;
    END
  END la_oenb[0]
  PIN la_oenb[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 672.610 0.000 672.890 4.000 ;
    END
  END la_oenb[100]
  PIN la_oenb[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 676.750 0.000 677.030 4.000 ;
    END
  END la_oenb[101]
  PIN la_oenb[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 680.890 0.000 681.170 4.000 ;
    END
  END la_oenb[102]
  PIN la_oenb[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 685.030 0.000 685.310 4.000 ;
    END
  END la_oenb[103]
  PIN la_oenb[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 689.170 0.000 689.450 4.000 ;
    END
  END la_oenb[104]
  PIN la_oenb[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 693.310 0.000 693.590 4.000 ;
    END
  END la_oenb[105]
  PIN la_oenb[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 697.450 0.000 697.730 4.000 ;
    END
  END la_oenb[106]
  PIN la_oenb[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 701.590 0.000 701.870 4.000 ;
    END
  END la_oenb[107]
  PIN la_oenb[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 705.730 0.000 706.010 4.000 ;
    END
  END la_oenb[108]
  PIN la_oenb[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 709.870 0.000 710.150 4.000 ;
    END
  END la_oenb[109]
  PIN la_oenb[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 300.010 0.000 300.290 4.000 ;
    END
  END la_oenb[10]
  PIN la_oenb[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 714.010 0.000 714.290 4.000 ;
    END
  END la_oenb[110]
  PIN la_oenb[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 718.150 0.000 718.430 4.000 ;
    END
  END la_oenb[111]
  PIN la_oenb[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 722.290 0.000 722.570 4.000 ;
    END
  END la_oenb[112]
  PIN la_oenb[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 726.430 0.000 726.710 4.000 ;
    END
  END la_oenb[113]
  PIN la_oenb[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 730.570 0.000 730.850 4.000 ;
    END
  END la_oenb[114]
  PIN la_oenb[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 734.710 0.000 734.990 4.000 ;
    END
  END la_oenb[115]
  PIN la_oenb[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 738.850 0.000 739.130 4.000 ;
    END
  END la_oenb[116]
  PIN la_oenb[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 742.990 0.000 743.270 4.000 ;
    END
  END la_oenb[117]
  PIN la_oenb[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 747.130 0.000 747.410 4.000 ;
    END
  END la_oenb[118]
  PIN la_oenb[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 751.270 0.000 751.550 4.000 ;
    END
  END la_oenb[119]
  PIN la_oenb[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 304.150 0.000 304.430 4.000 ;
    END
  END la_oenb[11]
  PIN la_oenb[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 755.410 0.000 755.690 4.000 ;
    END
  END la_oenb[120]
  PIN la_oenb[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 759.550 0.000 759.830 4.000 ;
    END
  END la_oenb[121]
  PIN la_oenb[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 763.690 0.000 763.970 4.000 ;
    END
  END la_oenb[122]
  PIN la_oenb[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 767.830 0.000 768.110 4.000 ;
    END
  END la_oenb[123]
  PIN la_oenb[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 771.970 0.000 772.250 4.000 ;
    END
  END la_oenb[124]
  PIN la_oenb[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 776.110 0.000 776.390 4.000 ;
    END
  END la_oenb[125]
  PIN la_oenb[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 780.250 0.000 780.530 4.000 ;
    END
  END la_oenb[126]
  PIN la_oenb[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 784.390 0.000 784.670 4.000 ;
    END
  END la_oenb[127]
  PIN la_oenb[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 308.290 0.000 308.570 4.000 ;
    END
  END la_oenb[12]
  PIN la_oenb[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 312.430 0.000 312.710 4.000 ;
    END
  END la_oenb[13]
  PIN la_oenb[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 316.570 0.000 316.850 4.000 ;
    END
  END la_oenb[14]
  PIN la_oenb[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 320.710 0.000 320.990 4.000 ;
    END
  END la_oenb[15]
  PIN la_oenb[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 324.850 0.000 325.130 4.000 ;
    END
  END la_oenb[16]
  PIN la_oenb[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 328.990 0.000 329.270 4.000 ;
    END
  END la_oenb[17]
  PIN la_oenb[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 333.130 0.000 333.410 4.000 ;
    END
  END la_oenb[18]
  PIN la_oenb[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 337.270 0.000 337.550 4.000 ;
    END
  END la_oenb[19]
  PIN la_oenb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 262.750 0.000 263.030 4.000 ;
    END
  END la_oenb[1]
  PIN la_oenb[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 341.410 0.000 341.690 4.000 ;
    END
  END la_oenb[20]
  PIN la_oenb[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 345.550 0.000 345.830 4.000 ;
    END
  END la_oenb[21]
  PIN la_oenb[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 349.690 0.000 349.970 4.000 ;
    END
  END la_oenb[22]
  PIN la_oenb[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 353.830 0.000 354.110 4.000 ;
    END
  END la_oenb[23]
  PIN la_oenb[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 357.970 0.000 358.250 4.000 ;
    END
  END la_oenb[24]
  PIN la_oenb[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 362.110 0.000 362.390 4.000 ;
    END
  END la_oenb[25]
  PIN la_oenb[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 366.250 0.000 366.530 4.000 ;
    END
  END la_oenb[26]
  PIN la_oenb[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 370.390 0.000 370.670 4.000 ;
    END
  END la_oenb[27]
  PIN la_oenb[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 374.530 0.000 374.810 4.000 ;
    END
  END la_oenb[28]
  PIN la_oenb[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 378.670 0.000 378.950 4.000 ;
    END
  END la_oenb[29]
  PIN la_oenb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 266.890 0.000 267.170 4.000 ;
    END
  END la_oenb[2]
  PIN la_oenb[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 382.810 0.000 383.090 4.000 ;
    END
  END la_oenb[30]
  PIN la_oenb[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 386.950 0.000 387.230 4.000 ;
    END
  END la_oenb[31]
  PIN la_oenb[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 391.090 0.000 391.370 4.000 ;
    END
  END la_oenb[32]
  PIN la_oenb[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 395.230 0.000 395.510 4.000 ;
    END
  END la_oenb[33]
  PIN la_oenb[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 399.370 0.000 399.650 4.000 ;
    END
  END la_oenb[34]
  PIN la_oenb[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 403.510 0.000 403.790 4.000 ;
    END
  END la_oenb[35]
  PIN la_oenb[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 407.650 0.000 407.930 4.000 ;
    END
  END la_oenb[36]
  PIN la_oenb[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 411.790 0.000 412.070 4.000 ;
    END
  END la_oenb[37]
  PIN la_oenb[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 415.930 0.000 416.210 4.000 ;
    END
  END la_oenb[38]
  PIN la_oenb[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 420.070 0.000 420.350 4.000 ;
    END
  END la_oenb[39]
  PIN la_oenb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 271.030 0.000 271.310 4.000 ;
    END
  END la_oenb[3]
  PIN la_oenb[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 424.210 0.000 424.490 4.000 ;
    END
  END la_oenb[40]
  PIN la_oenb[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 428.350 0.000 428.630 4.000 ;
    END
  END la_oenb[41]
  PIN la_oenb[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 432.490 0.000 432.770 4.000 ;
    END
  END la_oenb[42]
  PIN la_oenb[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 436.630 0.000 436.910 4.000 ;
    END
  END la_oenb[43]
  PIN la_oenb[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 440.770 0.000 441.050 4.000 ;
    END
  END la_oenb[44]
  PIN la_oenb[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 444.910 0.000 445.190 4.000 ;
    END
  END la_oenb[45]
  PIN la_oenb[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 449.050 0.000 449.330 4.000 ;
    END
  END la_oenb[46]
  PIN la_oenb[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 453.190 0.000 453.470 4.000 ;
    END
  END la_oenb[47]
  PIN la_oenb[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 457.330 0.000 457.610 4.000 ;
    END
  END la_oenb[48]
  PIN la_oenb[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 461.470 0.000 461.750 4.000 ;
    END
  END la_oenb[49]
  PIN la_oenb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 275.170 0.000 275.450 4.000 ;
    END
  END la_oenb[4]
  PIN la_oenb[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 465.610 0.000 465.890 4.000 ;
    END
  END la_oenb[50]
  PIN la_oenb[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 469.750 0.000 470.030 4.000 ;
    END
  END la_oenb[51]
  PIN la_oenb[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 473.890 0.000 474.170 4.000 ;
    END
  END la_oenb[52]
  PIN la_oenb[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 478.030 0.000 478.310 4.000 ;
    END
  END la_oenb[53]
  PIN la_oenb[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 482.170 0.000 482.450 4.000 ;
    END
  END la_oenb[54]
  PIN la_oenb[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 486.310 0.000 486.590 4.000 ;
    END
  END la_oenb[55]
  PIN la_oenb[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 490.450 0.000 490.730 4.000 ;
    END
  END la_oenb[56]
  PIN la_oenb[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 494.590 0.000 494.870 4.000 ;
    END
  END la_oenb[57]
  PIN la_oenb[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 498.730 0.000 499.010 4.000 ;
    END
  END la_oenb[58]
  PIN la_oenb[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 502.870 0.000 503.150 4.000 ;
    END
  END la_oenb[59]
  PIN la_oenb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 279.310 0.000 279.590 4.000 ;
    END
  END la_oenb[5]
  PIN la_oenb[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 507.010 0.000 507.290 4.000 ;
    END
  END la_oenb[60]
  PIN la_oenb[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 511.150 0.000 511.430 4.000 ;
    END
  END la_oenb[61]
  PIN la_oenb[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 515.290 0.000 515.570 4.000 ;
    END
  END la_oenb[62]
  PIN la_oenb[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 519.430 0.000 519.710 4.000 ;
    END
  END la_oenb[63]
  PIN la_oenb[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 523.570 0.000 523.850 4.000 ;
    END
  END la_oenb[64]
  PIN la_oenb[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 527.710 0.000 527.990 4.000 ;
    END
  END la_oenb[65]
  PIN la_oenb[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 531.850 0.000 532.130 4.000 ;
    END
  END la_oenb[66]
  PIN la_oenb[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 535.990 0.000 536.270 4.000 ;
    END
  END la_oenb[67]
  PIN la_oenb[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 540.130 0.000 540.410 4.000 ;
    END
  END la_oenb[68]
  PIN la_oenb[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 544.270 0.000 544.550 4.000 ;
    END
  END la_oenb[69]
  PIN la_oenb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 283.450 0.000 283.730 4.000 ;
    END
  END la_oenb[6]
  PIN la_oenb[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 548.410 0.000 548.690 4.000 ;
    END
  END la_oenb[70]
  PIN la_oenb[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 552.550 0.000 552.830 4.000 ;
    END
  END la_oenb[71]
  PIN la_oenb[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 556.690 0.000 556.970 4.000 ;
    END
  END la_oenb[72]
  PIN la_oenb[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 560.830 0.000 561.110 4.000 ;
    END
  END la_oenb[73]
  PIN la_oenb[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 564.970 0.000 565.250 4.000 ;
    END
  END la_oenb[74]
  PIN la_oenb[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 569.110 0.000 569.390 4.000 ;
    END
  END la_oenb[75]
  PIN la_oenb[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 573.250 0.000 573.530 4.000 ;
    END
  END la_oenb[76]
  PIN la_oenb[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 577.390 0.000 577.670 4.000 ;
    END
  END la_oenb[77]
  PIN la_oenb[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 581.530 0.000 581.810 4.000 ;
    END
  END la_oenb[78]
  PIN la_oenb[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 585.670 0.000 585.950 4.000 ;
    END
  END la_oenb[79]
  PIN la_oenb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 287.590 0.000 287.870 4.000 ;
    END
  END la_oenb[7]
  PIN la_oenb[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 589.810 0.000 590.090 4.000 ;
    END
  END la_oenb[80]
  PIN la_oenb[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 593.950 0.000 594.230 4.000 ;
    END
  END la_oenb[81]
  PIN la_oenb[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 598.090 0.000 598.370 4.000 ;
    END
  END la_oenb[82]
  PIN la_oenb[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 602.230 0.000 602.510 4.000 ;
    END
  END la_oenb[83]
  PIN la_oenb[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 606.370 0.000 606.650 4.000 ;
    END
  END la_oenb[84]
  PIN la_oenb[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 610.510 0.000 610.790 4.000 ;
    END
  END la_oenb[85]
  PIN la_oenb[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 614.650 0.000 614.930 4.000 ;
    END
  END la_oenb[86]
  PIN la_oenb[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 618.790 0.000 619.070 4.000 ;
    END
  END la_oenb[87]
  PIN la_oenb[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 622.930 0.000 623.210 4.000 ;
    END
  END la_oenb[88]
  PIN la_oenb[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 627.070 0.000 627.350 4.000 ;
    END
  END la_oenb[89]
  PIN la_oenb[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 291.730 0.000 292.010 4.000 ;
    END
  END la_oenb[8]
  PIN la_oenb[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 631.210 0.000 631.490 4.000 ;
    END
  END la_oenb[90]
  PIN la_oenb[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 635.350 0.000 635.630 4.000 ;
    END
  END la_oenb[91]
  PIN la_oenb[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 639.490 0.000 639.770 4.000 ;
    END
  END la_oenb[92]
  PIN la_oenb[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 643.630 0.000 643.910 4.000 ;
    END
  END la_oenb[93]
  PIN la_oenb[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 647.770 0.000 648.050 4.000 ;
    END
  END la_oenb[94]
  PIN la_oenb[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 651.910 0.000 652.190 4.000 ;
    END
  END la_oenb[95]
  PIN la_oenb[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 656.050 0.000 656.330 4.000 ;
    END
  END la_oenb[96]
  PIN la_oenb[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 660.190 0.000 660.470 4.000 ;
    END
  END la_oenb[97]
  PIN la_oenb[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 664.330 0.000 664.610 4.000 ;
    END
  END la_oenb[98]
  PIN la_oenb[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 668.470 0.000 668.750 4.000 ;
    END
  END la_oenb[99]
  PIN la_oenb[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 295.870 0.000 296.150 4.000 ;
    END
  END la_oenb[9]
  PIN user_clock2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 785.770 0.000 786.050 4.000 ;
    END
  END user_clock2
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 587.760 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 865.840 10.640 867.440 587.760 ;
    END
  END vssd1
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.570 0.000 109.850 4.000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 110.950 0.000 111.230 4.000 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.330 0.000 112.610 4.000 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 117.850 0.000 118.130 4.000 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 164.770 0.000 165.050 4.000 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 168.910 0.000 169.190 4.000 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.050 0.000 173.330 4.000 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 177.190 0.000 177.470 4.000 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 181.330 0.000 181.610 4.000 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 185.470 0.000 185.750 4.000 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 189.610 0.000 189.890 4.000 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 193.750 0.000 194.030 4.000 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 197.890 0.000 198.170 4.000 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.030 0.000 202.310 4.000 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 123.370 0.000 123.650 4.000 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 206.170 0.000 206.450 4.000 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 210.310 0.000 210.590 4.000 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 214.450 0.000 214.730 4.000 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 218.590 0.000 218.870 4.000 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 222.730 0.000 223.010 4.000 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 226.870 0.000 227.150 4.000 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 231.010 0.000 231.290 4.000 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 235.150 0.000 235.430 4.000 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 239.290 0.000 239.570 4.000 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 243.430 0.000 243.710 4.000 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.890 0.000 129.170 4.000 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 247.570 0.000 247.850 4.000 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 251.710 0.000 251.990 4.000 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 134.410 0.000 134.690 4.000 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 139.930 0.000 140.210 4.000 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.070 0.000 144.350 4.000 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 148.210 0.000 148.490 4.000 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 152.350 0.000 152.630 4.000 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 156.490 0.000 156.770 4.000 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 160.630 0.000 160.910 4.000 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 113.710 0.000 113.990 4.000 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.230 0.000 119.510 4.000 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 166.150 0.000 166.430 4.000 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 170.290 0.000 170.570 4.000 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 174.430 0.000 174.710 4.000 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 178.570 0.000 178.850 4.000 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 182.710 0.000 182.990 4.000 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 186.850 0.000 187.130 4.000 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.990 0.000 191.270 4.000 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 195.130 0.000 195.410 4.000 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 199.270 0.000 199.550 4.000 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 203.410 0.000 203.690 4.000 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 124.750 0.000 125.030 4.000 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 207.550 0.000 207.830 4.000 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 211.690 0.000 211.970 4.000 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 215.830 0.000 216.110 4.000 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 219.970 0.000 220.250 4.000 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 224.110 0.000 224.390 4.000 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 228.250 0.000 228.530 4.000 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 232.390 0.000 232.670 4.000 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 236.530 0.000 236.810 4.000 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 240.670 0.000 240.950 4.000 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 244.810 0.000 245.090 4.000 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 130.270 0.000 130.550 4.000 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 248.950 0.000 249.230 4.000 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 253.090 0.000 253.370 4.000 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.790 0.000 136.070 4.000 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 141.310 0.000 141.590 4.000 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 145.450 0.000 145.730 4.000 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 149.590 0.000 149.870 4.000 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 153.730 0.000 154.010 4.000 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.870 0.000 158.150 4.000 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 162.010 0.000 162.290 4.000 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 120.610 0.000 120.890 4.000 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.530 0.000 167.810 4.000 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 171.670 0.000 171.950 4.000 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 175.810 0.000 176.090 4.000 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 179.950 0.000 180.230 4.000 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 184.090 0.000 184.370 4.000 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 188.230 0.000 188.510 4.000 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 192.370 0.000 192.650 4.000 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.510 0.000 196.790 4.000 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 200.650 0.000 200.930 4.000 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 204.790 0.000 205.070 4.000 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 126.130 0.000 126.410 4.000 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.930 0.000 209.210 4.000 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 213.070 0.000 213.350 4.000 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 217.210 0.000 217.490 4.000 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 221.350 0.000 221.630 4.000 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 225.490 0.000 225.770 4.000 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 229.630 0.000 229.910 4.000 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 233.770 0.000 234.050 4.000 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 237.910 0.000 238.190 4.000 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 242.050 0.000 242.330 4.000 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 246.190 0.000 246.470 4.000 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 131.650 0.000 131.930 4.000 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 250.330 0.000 250.610 4.000 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 254.470 0.000 254.750 4.000 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 137.170 0.000 137.450 4.000 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 142.690 0.000 142.970 4.000 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 146.830 0.000 147.110 4.000 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.970 0.000 151.250 4.000 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 155.110 0.000 155.390 4.000 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 159.250 0.000 159.530 4.000 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 163.390 0.000 163.670 4.000 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.990 0.000 122.270 4.000 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 127.510 0.000 127.790 4.000 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 133.030 0.000 133.310 4.000 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.550 0.000 138.830 4.000 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 115.090 0.000 115.370 4.000 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.470 0.000 116.750 4.000 ;
    END
  END wbs_we_i
  OBS
      LAYER nwell ;
        RECT 5.330 583.385 894.430 586.215 ;
        RECT 5.330 577.945 894.430 580.775 ;
        RECT 5.330 572.505 894.430 575.335 ;
        RECT 5.330 567.065 894.430 569.895 ;
        RECT 5.330 561.625 894.430 564.455 ;
        RECT 5.330 556.185 894.430 559.015 ;
        RECT 5.330 550.745 894.430 553.575 ;
        RECT 5.330 545.305 894.430 548.135 ;
        RECT 5.330 539.865 894.430 542.695 ;
        RECT 5.330 534.425 894.430 537.255 ;
        RECT 5.330 528.985 894.430 531.815 ;
        RECT 5.330 523.545 894.430 526.375 ;
        RECT 5.330 518.105 894.430 520.935 ;
        RECT 5.330 512.665 894.430 515.495 ;
        RECT 5.330 507.225 894.430 510.055 ;
        RECT 5.330 501.785 894.430 504.615 ;
        RECT 5.330 496.345 894.430 499.175 ;
        RECT 5.330 490.905 894.430 493.735 ;
        RECT 5.330 485.465 894.430 488.295 ;
        RECT 5.330 480.025 894.430 482.855 ;
        RECT 5.330 474.585 894.430 477.415 ;
        RECT 5.330 469.145 894.430 471.975 ;
        RECT 5.330 463.705 894.430 466.535 ;
        RECT 5.330 458.265 894.430 461.095 ;
        RECT 5.330 452.825 894.430 455.655 ;
        RECT 5.330 447.385 894.430 450.215 ;
        RECT 5.330 441.945 894.430 444.775 ;
        RECT 5.330 436.505 894.430 439.335 ;
        RECT 5.330 431.065 894.430 433.895 ;
        RECT 5.330 425.625 894.430 428.455 ;
        RECT 5.330 420.185 894.430 423.015 ;
        RECT 5.330 414.745 894.430 417.575 ;
        RECT 5.330 409.305 894.430 412.135 ;
        RECT 5.330 403.865 894.430 406.695 ;
        RECT 5.330 398.425 894.430 401.255 ;
        RECT 5.330 392.985 894.430 395.815 ;
        RECT 5.330 387.545 894.430 390.375 ;
        RECT 5.330 382.105 894.430 384.935 ;
        RECT 5.330 376.665 894.430 379.495 ;
        RECT 5.330 371.225 894.430 374.055 ;
        RECT 5.330 365.785 894.430 368.615 ;
        RECT 5.330 360.345 894.430 363.175 ;
        RECT 5.330 354.905 894.430 357.735 ;
        RECT 5.330 349.465 894.430 352.295 ;
        RECT 5.330 344.025 894.430 346.855 ;
        RECT 5.330 338.585 894.430 341.415 ;
        RECT 5.330 333.145 894.430 335.975 ;
        RECT 5.330 327.705 894.430 330.535 ;
        RECT 5.330 322.265 894.430 325.095 ;
        RECT 5.330 316.825 894.430 319.655 ;
        RECT 5.330 311.385 894.430 314.215 ;
        RECT 5.330 305.945 894.430 308.775 ;
        RECT 5.330 300.505 894.430 303.335 ;
        RECT 5.330 295.065 894.430 297.895 ;
        RECT 5.330 289.625 894.430 292.455 ;
        RECT 5.330 284.185 894.430 287.015 ;
        RECT 5.330 278.745 894.430 281.575 ;
        RECT 5.330 273.305 894.430 276.135 ;
        RECT 5.330 267.865 894.430 270.695 ;
        RECT 5.330 262.425 894.430 265.255 ;
        RECT 5.330 256.985 894.430 259.815 ;
        RECT 5.330 251.545 894.430 254.375 ;
        RECT 5.330 246.105 894.430 248.935 ;
        RECT 5.330 240.665 894.430 243.495 ;
        RECT 5.330 235.225 894.430 238.055 ;
        RECT 5.330 229.785 894.430 232.615 ;
        RECT 5.330 224.345 894.430 227.175 ;
        RECT 5.330 218.905 894.430 221.735 ;
        RECT 5.330 213.465 894.430 216.295 ;
        RECT 5.330 208.025 894.430 210.855 ;
        RECT 5.330 202.585 894.430 205.415 ;
        RECT 5.330 197.145 894.430 199.975 ;
        RECT 5.330 191.705 894.430 194.535 ;
        RECT 5.330 186.265 894.430 189.095 ;
        RECT 5.330 180.825 894.430 183.655 ;
        RECT 5.330 175.385 894.430 178.215 ;
        RECT 5.330 169.945 894.430 172.775 ;
        RECT 5.330 164.505 894.430 167.335 ;
        RECT 5.330 159.065 894.430 161.895 ;
        RECT 5.330 153.625 894.430 156.455 ;
        RECT 5.330 148.185 894.430 151.015 ;
        RECT 5.330 142.745 894.430 145.575 ;
        RECT 5.330 137.305 894.430 140.135 ;
        RECT 5.330 131.865 894.430 134.695 ;
        RECT 5.330 126.425 894.430 129.255 ;
        RECT 5.330 120.985 894.430 123.815 ;
        RECT 5.330 115.545 894.430 118.375 ;
        RECT 5.330 110.105 894.430 112.935 ;
        RECT 5.330 104.665 894.430 107.495 ;
        RECT 5.330 99.225 894.430 102.055 ;
        RECT 5.330 93.785 894.430 96.615 ;
        RECT 5.330 88.345 894.430 91.175 ;
        RECT 5.330 82.905 894.430 85.735 ;
        RECT 5.330 77.465 894.430 80.295 ;
        RECT 5.330 72.025 894.430 74.855 ;
        RECT 5.330 66.585 894.430 69.415 ;
        RECT 5.330 61.145 894.430 63.975 ;
        RECT 5.330 55.705 894.430 58.535 ;
        RECT 5.330 50.265 894.430 53.095 ;
        RECT 5.330 44.825 894.430 47.655 ;
        RECT 5.330 39.385 894.430 42.215 ;
        RECT 5.330 33.945 894.430 36.775 ;
        RECT 5.330 28.505 894.430 31.335 ;
        RECT 5.330 23.065 894.430 25.895 ;
        RECT 5.330 17.625 894.430 20.455 ;
        RECT 5.330 12.185 894.430 15.015 ;
      LAYER li1 ;
        RECT 5.520 10.795 894.240 587.605 ;
      LAYER met1 ;
        RECT 5.520 3.100 894.240 587.760 ;
      LAYER met2 ;
        RECT 16.290 595.720 23.270 596.770 ;
        RECT 24.110 595.720 31.090 596.770 ;
        RECT 31.930 595.720 38.910 596.770 ;
        RECT 39.750 595.720 46.730 596.770 ;
        RECT 47.570 595.720 54.550 596.770 ;
        RECT 55.390 595.720 62.370 596.770 ;
        RECT 63.210 595.720 70.190 596.770 ;
        RECT 71.030 595.720 78.010 596.770 ;
        RECT 78.850 595.720 85.830 596.770 ;
        RECT 86.670 595.720 93.650 596.770 ;
        RECT 94.490 595.720 101.470 596.770 ;
        RECT 102.310 595.720 109.290 596.770 ;
        RECT 110.130 595.720 117.110 596.770 ;
        RECT 117.950 595.720 124.930 596.770 ;
        RECT 125.770 595.720 132.750 596.770 ;
        RECT 133.590 595.720 140.570 596.770 ;
        RECT 141.410 595.720 148.390 596.770 ;
        RECT 149.230 595.720 156.210 596.770 ;
        RECT 157.050 595.720 164.030 596.770 ;
        RECT 164.870 595.720 171.850 596.770 ;
        RECT 172.690 595.720 179.670 596.770 ;
        RECT 180.510 595.720 187.490 596.770 ;
        RECT 188.330 595.720 195.310 596.770 ;
        RECT 196.150 595.720 203.130 596.770 ;
        RECT 203.970 595.720 210.950 596.770 ;
        RECT 211.790 595.720 218.770 596.770 ;
        RECT 219.610 595.720 226.590 596.770 ;
        RECT 227.430 595.720 234.410 596.770 ;
        RECT 235.250 595.720 242.230 596.770 ;
        RECT 243.070 595.720 250.050 596.770 ;
        RECT 250.890 595.720 257.870 596.770 ;
        RECT 258.710 595.720 265.690 596.770 ;
        RECT 266.530 595.720 273.510 596.770 ;
        RECT 274.350 595.720 281.330 596.770 ;
        RECT 282.170 595.720 289.150 596.770 ;
        RECT 289.990 595.720 296.970 596.770 ;
        RECT 297.810 595.720 304.790 596.770 ;
        RECT 305.630 595.720 312.610 596.770 ;
        RECT 313.450 595.720 320.430 596.770 ;
        RECT 321.270 595.720 328.250 596.770 ;
        RECT 329.090 595.720 336.070 596.770 ;
        RECT 336.910 595.720 343.890 596.770 ;
        RECT 344.730 595.720 351.710 596.770 ;
        RECT 352.550 595.720 359.530 596.770 ;
        RECT 360.370 595.720 367.350 596.770 ;
        RECT 368.190 595.720 375.170 596.770 ;
        RECT 376.010 595.720 382.990 596.770 ;
        RECT 383.830 595.720 390.810 596.770 ;
        RECT 391.650 595.720 398.630 596.770 ;
        RECT 399.470 595.720 406.450 596.770 ;
        RECT 407.290 595.720 414.270 596.770 ;
        RECT 415.110 595.720 422.090 596.770 ;
        RECT 422.930 595.720 429.910 596.770 ;
        RECT 430.750 595.720 437.730 596.770 ;
        RECT 438.570 595.720 445.550 596.770 ;
        RECT 446.390 595.720 453.370 596.770 ;
        RECT 454.210 595.720 461.190 596.770 ;
        RECT 462.030 595.720 469.010 596.770 ;
        RECT 469.850 595.720 476.830 596.770 ;
        RECT 477.670 595.720 484.650 596.770 ;
        RECT 485.490 595.720 492.470 596.770 ;
        RECT 493.310 595.720 500.290 596.770 ;
        RECT 501.130 595.720 508.110 596.770 ;
        RECT 508.950 595.720 515.930 596.770 ;
        RECT 516.770 595.720 523.750 596.770 ;
        RECT 524.590 595.720 531.570 596.770 ;
        RECT 532.410 595.720 539.390 596.770 ;
        RECT 540.230 595.720 547.210 596.770 ;
        RECT 548.050 595.720 555.030 596.770 ;
        RECT 555.870 595.720 562.850 596.770 ;
        RECT 563.690 595.720 570.670 596.770 ;
        RECT 571.510 595.720 578.490 596.770 ;
        RECT 579.330 595.720 586.310 596.770 ;
        RECT 587.150 595.720 594.130 596.770 ;
        RECT 594.970 595.720 601.950 596.770 ;
        RECT 602.790 595.720 609.770 596.770 ;
        RECT 610.610 595.720 617.590 596.770 ;
        RECT 618.430 595.720 625.410 596.770 ;
        RECT 626.250 595.720 633.230 596.770 ;
        RECT 634.070 595.720 641.050 596.770 ;
        RECT 641.890 595.720 648.870 596.770 ;
        RECT 649.710 595.720 656.690 596.770 ;
        RECT 657.530 595.720 664.510 596.770 ;
        RECT 665.350 595.720 672.330 596.770 ;
        RECT 673.170 595.720 680.150 596.770 ;
        RECT 680.990 595.720 687.970 596.770 ;
        RECT 688.810 595.720 695.790 596.770 ;
        RECT 696.630 595.720 703.610 596.770 ;
        RECT 704.450 595.720 711.430 596.770 ;
        RECT 712.270 595.720 719.250 596.770 ;
        RECT 720.090 595.720 727.070 596.770 ;
        RECT 727.910 595.720 734.890 596.770 ;
        RECT 735.730 595.720 742.710 596.770 ;
        RECT 743.550 595.720 750.530 596.770 ;
        RECT 751.370 595.720 758.350 596.770 ;
        RECT 759.190 595.720 766.170 596.770 ;
        RECT 767.010 595.720 773.990 596.770 ;
        RECT 774.830 595.720 781.810 596.770 ;
        RECT 782.650 595.720 789.630 596.770 ;
        RECT 790.470 595.720 797.450 596.770 ;
        RECT 798.290 595.720 805.270 596.770 ;
        RECT 806.110 595.720 813.090 596.770 ;
        RECT 813.930 595.720 820.910 596.770 ;
        RECT 821.750 595.720 828.730 596.770 ;
        RECT 829.570 595.720 836.550 596.770 ;
        RECT 837.390 595.720 844.370 596.770 ;
        RECT 845.210 595.720 852.190 596.770 ;
        RECT 853.030 595.720 860.010 596.770 ;
        RECT 860.850 595.720 867.830 596.770 ;
        RECT 868.670 595.720 875.650 596.770 ;
        RECT 876.490 595.720 883.470 596.770 ;
        RECT 884.310 595.720 891.290 596.770 ;
        RECT 16.010 4.280 891.840 595.720 ;
        RECT 16.010 3.070 109.290 4.280 ;
        RECT 110.130 3.070 110.670 4.280 ;
        RECT 111.510 3.070 112.050 4.280 ;
        RECT 112.890 3.070 113.430 4.280 ;
        RECT 114.270 3.070 114.810 4.280 ;
        RECT 115.650 3.070 116.190 4.280 ;
        RECT 117.030 3.070 117.570 4.280 ;
        RECT 118.410 3.070 118.950 4.280 ;
        RECT 119.790 3.070 120.330 4.280 ;
        RECT 121.170 3.070 121.710 4.280 ;
        RECT 122.550 3.070 123.090 4.280 ;
        RECT 123.930 3.070 124.470 4.280 ;
        RECT 125.310 3.070 125.850 4.280 ;
        RECT 126.690 3.070 127.230 4.280 ;
        RECT 128.070 3.070 128.610 4.280 ;
        RECT 129.450 3.070 129.990 4.280 ;
        RECT 130.830 3.070 131.370 4.280 ;
        RECT 132.210 3.070 132.750 4.280 ;
        RECT 133.590 3.070 134.130 4.280 ;
        RECT 134.970 3.070 135.510 4.280 ;
        RECT 136.350 3.070 136.890 4.280 ;
        RECT 137.730 3.070 138.270 4.280 ;
        RECT 139.110 3.070 139.650 4.280 ;
        RECT 140.490 3.070 141.030 4.280 ;
        RECT 141.870 3.070 142.410 4.280 ;
        RECT 143.250 3.070 143.790 4.280 ;
        RECT 144.630 3.070 145.170 4.280 ;
        RECT 146.010 3.070 146.550 4.280 ;
        RECT 147.390 3.070 147.930 4.280 ;
        RECT 148.770 3.070 149.310 4.280 ;
        RECT 150.150 3.070 150.690 4.280 ;
        RECT 151.530 3.070 152.070 4.280 ;
        RECT 152.910 3.070 153.450 4.280 ;
        RECT 154.290 3.070 154.830 4.280 ;
        RECT 155.670 3.070 156.210 4.280 ;
        RECT 157.050 3.070 157.590 4.280 ;
        RECT 158.430 3.070 158.970 4.280 ;
        RECT 159.810 3.070 160.350 4.280 ;
        RECT 161.190 3.070 161.730 4.280 ;
        RECT 162.570 3.070 163.110 4.280 ;
        RECT 163.950 3.070 164.490 4.280 ;
        RECT 165.330 3.070 165.870 4.280 ;
        RECT 166.710 3.070 167.250 4.280 ;
        RECT 168.090 3.070 168.630 4.280 ;
        RECT 169.470 3.070 170.010 4.280 ;
        RECT 170.850 3.070 171.390 4.280 ;
        RECT 172.230 3.070 172.770 4.280 ;
        RECT 173.610 3.070 174.150 4.280 ;
        RECT 174.990 3.070 175.530 4.280 ;
        RECT 176.370 3.070 176.910 4.280 ;
        RECT 177.750 3.070 178.290 4.280 ;
        RECT 179.130 3.070 179.670 4.280 ;
        RECT 180.510 3.070 181.050 4.280 ;
        RECT 181.890 3.070 182.430 4.280 ;
        RECT 183.270 3.070 183.810 4.280 ;
        RECT 184.650 3.070 185.190 4.280 ;
        RECT 186.030 3.070 186.570 4.280 ;
        RECT 187.410 3.070 187.950 4.280 ;
        RECT 188.790 3.070 189.330 4.280 ;
        RECT 190.170 3.070 190.710 4.280 ;
        RECT 191.550 3.070 192.090 4.280 ;
        RECT 192.930 3.070 193.470 4.280 ;
        RECT 194.310 3.070 194.850 4.280 ;
        RECT 195.690 3.070 196.230 4.280 ;
        RECT 197.070 3.070 197.610 4.280 ;
        RECT 198.450 3.070 198.990 4.280 ;
        RECT 199.830 3.070 200.370 4.280 ;
        RECT 201.210 3.070 201.750 4.280 ;
        RECT 202.590 3.070 203.130 4.280 ;
        RECT 203.970 3.070 204.510 4.280 ;
        RECT 205.350 3.070 205.890 4.280 ;
        RECT 206.730 3.070 207.270 4.280 ;
        RECT 208.110 3.070 208.650 4.280 ;
        RECT 209.490 3.070 210.030 4.280 ;
        RECT 210.870 3.070 211.410 4.280 ;
        RECT 212.250 3.070 212.790 4.280 ;
        RECT 213.630 3.070 214.170 4.280 ;
        RECT 215.010 3.070 215.550 4.280 ;
        RECT 216.390 3.070 216.930 4.280 ;
        RECT 217.770 3.070 218.310 4.280 ;
        RECT 219.150 3.070 219.690 4.280 ;
        RECT 220.530 3.070 221.070 4.280 ;
        RECT 221.910 3.070 222.450 4.280 ;
        RECT 223.290 3.070 223.830 4.280 ;
        RECT 224.670 3.070 225.210 4.280 ;
        RECT 226.050 3.070 226.590 4.280 ;
        RECT 227.430 3.070 227.970 4.280 ;
        RECT 228.810 3.070 229.350 4.280 ;
        RECT 230.190 3.070 230.730 4.280 ;
        RECT 231.570 3.070 232.110 4.280 ;
        RECT 232.950 3.070 233.490 4.280 ;
        RECT 234.330 3.070 234.870 4.280 ;
        RECT 235.710 3.070 236.250 4.280 ;
        RECT 237.090 3.070 237.630 4.280 ;
        RECT 238.470 3.070 239.010 4.280 ;
        RECT 239.850 3.070 240.390 4.280 ;
        RECT 241.230 3.070 241.770 4.280 ;
        RECT 242.610 3.070 243.150 4.280 ;
        RECT 243.990 3.070 244.530 4.280 ;
        RECT 245.370 3.070 245.910 4.280 ;
        RECT 246.750 3.070 247.290 4.280 ;
        RECT 248.130 3.070 248.670 4.280 ;
        RECT 249.510 3.070 250.050 4.280 ;
        RECT 250.890 3.070 251.430 4.280 ;
        RECT 252.270 3.070 252.810 4.280 ;
        RECT 253.650 3.070 254.190 4.280 ;
        RECT 255.030 3.070 255.570 4.280 ;
        RECT 256.410 3.070 256.950 4.280 ;
        RECT 257.790 3.070 258.330 4.280 ;
        RECT 259.170 3.070 259.710 4.280 ;
        RECT 260.550 3.070 261.090 4.280 ;
        RECT 261.930 3.070 262.470 4.280 ;
        RECT 263.310 3.070 263.850 4.280 ;
        RECT 264.690 3.070 265.230 4.280 ;
        RECT 266.070 3.070 266.610 4.280 ;
        RECT 267.450 3.070 267.990 4.280 ;
        RECT 268.830 3.070 269.370 4.280 ;
        RECT 270.210 3.070 270.750 4.280 ;
        RECT 271.590 3.070 272.130 4.280 ;
        RECT 272.970 3.070 273.510 4.280 ;
        RECT 274.350 3.070 274.890 4.280 ;
        RECT 275.730 3.070 276.270 4.280 ;
        RECT 277.110 3.070 277.650 4.280 ;
        RECT 278.490 3.070 279.030 4.280 ;
        RECT 279.870 3.070 280.410 4.280 ;
        RECT 281.250 3.070 281.790 4.280 ;
        RECT 282.630 3.070 283.170 4.280 ;
        RECT 284.010 3.070 284.550 4.280 ;
        RECT 285.390 3.070 285.930 4.280 ;
        RECT 286.770 3.070 287.310 4.280 ;
        RECT 288.150 3.070 288.690 4.280 ;
        RECT 289.530 3.070 290.070 4.280 ;
        RECT 290.910 3.070 291.450 4.280 ;
        RECT 292.290 3.070 292.830 4.280 ;
        RECT 293.670 3.070 294.210 4.280 ;
        RECT 295.050 3.070 295.590 4.280 ;
        RECT 296.430 3.070 296.970 4.280 ;
        RECT 297.810 3.070 298.350 4.280 ;
        RECT 299.190 3.070 299.730 4.280 ;
        RECT 300.570 3.070 301.110 4.280 ;
        RECT 301.950 3.070 302.490 4.280 ;
        RECT 303.330 3.070 303.870 4.280 ;
        RECT 304.710 3.070 305.250 4.280 ;
        RECT 306.090 3.070 306.630 4.280 ;
        RECT 307.470 3.070 308.010 4.280 ;
        RECT 308.850 3.070 309.390 4.280 ;
        RECT 310.230 3.070 310.770 4.280 ;
        RECT 311.610 3.070 312.150 4.280 ;
        RECT 312.990 3.070 313.530 4.280 ;
        RECT 314.370 3.070 314.910 4.280 ;
        RECT 315.750 3.070 316.290 4.280 ;
        RECT 317.130 3.070 317.670 4.280 ;
        RECT 318.510 3.070 319.050 4.280 ;
        RECT 319.890 3.070 320.430 4.280 ;
        RECT 321.270 3.070 321.810 4.280 ;
        RECT 322.650 3.070 323.190 4.280 ;
        RECT 324.030 3.070 324.570 4.280 ;
        RECT 325.410 3.070 325.950 4.280 ;
        RECT 326.790 3.070 327.330 4.280 ;
        RECT 328.170 3.070 328.710 4.280 ;
        RECT 329.550 3.070 330.090 4.280 ;
        RECT 330.930 3.070 331.470 4.280 ;
        RECT 332.310 3.070 332.850 4.280 ;
        RECT 333.690 3.070 334.230 4.280 ;
        RECT 335.070 3.070 335.610 4.280 ;
        RECT 336.450 3.070 336.990 4.280 ;
        RECT 337.830 3.070 338.370 4.280 ;
        RECT 339.210 3.070 339.750 4.280 ;
        RECT 340.590 3.070 341.130 4.280 ;
        RECT 341.970 3.070 342.510 4.280 ;
        RECT 343.350 3.070 343.890 4.280 ;
        RECT 344.730 3.070 345.270 4.280 ;
        RECT 346.110 3.070 346.650 4.280 ;
        RECT 347.490 3.070 348.030 4.280 ;
        RECT 348.870 3.070 349.410 4.280 ;
        RECT 350.250 3.070 350.790 4.280 ;
        RECT 351.630 3.070 352.170 4.280 ;
        RECT 353.010 3.070 353.550 4.280 ;
        RECT 354.390 3.070 354.930 4.280 ;
        RECT 355.770 3.070 356.310 4.280 ;
        RECT 357.150 3.070 357.690 4.280 ;
        RECT 358.530 3.070 359.070 4.280 ;
        RECT 359.910 3.070 360.450 4.280 ;
        RECT 361.290 3.070 361.830 4.280 ;
        RECT 362.670 3.070 363.210 4.280 ;
        RECT 364.050 3.070 364.590 4.280 ;
        RECT 365.430 3.070 365.970 4.280 ;
        RECT 366.810 3.070 367.350 4.280 ;
        RECT 368.190 3.070 368.730 4.280 ;
        RECT 369.570 3.070 370.110 4.280 ;
        RECT 370.950 3.070 371.490 4.280 ;
        RECT 372.330 3.070 372.870 4.280 ;
        RECT 373.710 3.070 374.250 4.280 ;
        RECT 375.090 3.070 375.630 4.280 ;
        RECT 376.470 3.070 377.010 4.280 ;
        RECT 377.850 3.070 378.390 4.280 ;
        RECT 379.230 3.070 379.770 4.280 ;
        RECT 380.610 3.070 381.150 4.280 ;
        RECT 381.990 3.070 382.530 4.280 ;
        RECT 383.370 3.070 383.910 4.280 ;
        RECT 384.750 3.070 385.290 4.280 ;
        RECT 386.130 3.070 386.670 4.280 ;
        RECT 387.510 3.070 388.050 4.280 ;
        RECT 388.890 3.070 389.430 4.280 ;
        RECT 390.270 3.070 390.810 4.280 ;
        RECT 391.650 3.070 392.190 4.280 ;
        RECT 393.030 3.070 393.570 4.280 ;
        RECT 394.410 3.070 394.950 4.280 ;
        RECT 395.790 3.070 396.330 4.280 ;
        RECT 397.170 3.070 397.710 4.280 ;
        RECT 398.550 3.070 399.090 4.280 ;
        RECT 399.930 3.070 400.470 4.280 ;
        RECT 401.310 3.070 401.850 4.280 ;
        RECT 402.690 3.070 403.230 4.280 ;
        RECT 404.070 3.070 404.610 4.280 ;
        RECT 405.450 3.070 405.990 4.280 ;
        RECT 406.830 3.070 407.370 4.280 ;
        RECT 408.210 3.070 408.750 4.280 ;
        RECT 409.590 3.070 410.130 4.280 ;
        RECT 410.970 3.070 411.510 4.280 ;
        RECT 412.350 3.070 412.890 4.280 ;
        RECT 413.730 3.070 414.270 4.280 ;
        RECT 415.110 3.070 415.650 4.280 ;
        RECT 416.490 3.070 417.030 4.280 ;
        RECT 417.870 3.070 418.410 4.280 ;
        RECT 419.250 3.070 419.790 4.280 ;
        RECT 420.630 3.070 421.170 4.280 ;
        RECT 422.010 3.070 422.550 4.280 ;
        RECT 423.390 3.070 423.930 4.280 ;
        RECT 424.770 3.070 425.310 4.280 ;
        RECT 426.150 3.070 426.690 4.280 ;
        RECT 427.530 3.070 428.070 4.280 ;
        RECT 428.910 3.070 429.450 4.280 ;
        RECT 430.290 3.070 430.830 4.280 ;
        RECT 431.670 3.070 432.210 4.280 ;
        RECT 433.050 3.070 433.590 4.280 ;
        RECT 434.430 3.070 434.970 4.280 ;
        RECT 435.810 3.070 436.350 4.280 ;
        RECT 437.190 3.070 437.730 4.280 ;
        RECT 438.570 3.070 439.110 4.280 ;
        RECT 439.950 3.070 440.490 4.280 ;
        RECT 441.330 3.070 441.870 4.280 ;
        RECT 442.710 3.070 443.250 4.280 ;
        RECT 444.090 3.070 444.630 4.280 ;
        RECT 445.470 3.070 446.010 4.280 ;
        RECT 446.850 3.070 447.390 4.280 ;
        RECT 448.230 3.070 448.770 4.280 ;
        RECT 449.610 3.070 450.150 4.280 ;
        RECT 450.990 3.070 451.530 4.280 ;
        RECT 452.370 3.070 452.910 4.280 ;
        RECT 453.750 3.070 454.290 4.280 ;
        RECT 455.130 3.070 455.670 4.280 ;
        RECT 456.510 3.070 457.050 4.280 ;
        RECT 457.890 3.070 458.430 4.280 ;
        RECT 459.270 3.070 459.810 4.280 ;
        RECT 460.650 3.070 461.190 4.280 ;
        RECT 462.030 3.070 462.570 4.280 ;
        RECT 463.410 3.070 463.950 4.280 ;
        RECT 464.790 3.070 465.330 4.280 ;
        RECT 466.170 3.070 466.710 4.280 ;
        RECT 467.550 3.070 468.090 4.280 ;
        RECT 468.930 3.070 469.470 4.280 ;
        RECT 470.310 3.070 470.850 4.280 ;
        RECT 471.690 3.070 472.230 4.280 ;
        RECT 473.070 3.070 473.610 4.280 ;
        RECT 474.450 3.070 474.990 4.280 ;
        RECT 475.830 3.070 476.370 4.280 ;
        RECT 477.210 3.070 477.750 4.280 ;
        RECT 478.590 3.070 479.130 4.280 ;
        RECT 479.970 3.070 480.510 4.280 ;
        RECT 481.350 3.070 481.890 4.280 ;
        RECT 482.730 3.070 483.270 4.280 ;
        RECT 484.110 3.070 484.650 4.280 ;
        RECT 485.490 3.070 486.030 4.280 ;
        RECT 486.870 3.070 487.410 4.280 ;
        RECT 488.250 3.070 488.790 4.280 ;
        RECT 489.630 3.070 490.170 4.280 ;
        RECT 491.010 3.070 491.550 4.280 ;
        RECT 492.390 3.070 492.930 4.280 ;
        RECT 493.770 3.070 494.310 4.280 ;
        RECT 495.150 3.070 495.690 4.280 ;
        RECT 496.530 3.070 497.070 4.280 ;
        RECT 497.910 3.070 498.450 4.280 ;
        RECT 499.290 3.070 499.830 4.280 ;
        RECT 500.670 3.070 501.210 4.280 ;
        RECT 502.050 3.070 502.590 4.280 ;
        RECT 503.430 3.070 503.970 4.280 ;
        RECT 504.810 3.070 505.350 4.280 ;
        RECT 506.190 3.070 506.730 4.280 ;
        RECT 507.570 3.070 508.110 4.280 ;
        RECT 508.950 3.070 509.490 4.280 ;
        RECT 510.330 3.070 510.870 4.280 ;
        RECT 511.710 3.070 512.250 4.280 ;
        RECT 513.090 3.070 513.630 4.280 ;
        RECT 514.470 3.070 515.010 4.280 ;
        RECT 515.850 3.070 516.390 4.280 ;
        RECT 517.230 3.070 517.770 4.280 ;
        RECT 518.610 3.070 519.150 4.280 ;
        RECT 519.990 3.070 520.530 4.280 ;
        RECT 521.370 3.070 521.910 4.280 ;
        RECT 522.750 3.070 523.290 4.280 ;
        RECT 524.130 3.070 524.670 4.280 ;
        RECT 525.510 3.070 526.050 4.280 ;
        RECT 526.890 3.070 527.430 4.280 ;
        RECT 528.270 3.070 528.810 4.280 ;
        RECT 529.650 3.070 530.190 4.280 ;
        RECT 531.030 3.070 531.570 4.280 ;
        RECT 532.410 3.070 532.950 4.280 ;
        RECT 533.790 3.070 534.330 4.280 ;
        RECT 535.170 3.070 535.710 4.280 ;
        RECT 536.550 3.070 537.090 4.280 ;
        RECT 537.930 3.070 538.470 4.280 ;
        RECT 539.310 3.070 539.850 4.280 ;
        RECT 540.690 3.070 541.230 4.280 ;
        RECT 542.070 3.070 542.610 4.280 ;
        RECT 543.450 3.070 543.990 4.280 ;
        RECT 544.830 3.070 545.370 4.280 ;
        RECT 546.210 3.070 546.750 4.280 ;
        RECT 547.590 3.070 548.130 4.280 ;
        RECT 548.970 3.070 549.510 4.280 ;
        RECT 550.350 3.070 550.890 4.280 ;
        RECT 551.730 3.070 552.270 4.280 ;
        RECT 553.110 3.070 553.650 4.280 ;
        RECT 554.490 3.070 555.030 4.280 ;
        RECT 555.870 3.070 556.410 4.280 ;
        RECT 557.250 3.070 557.790 4.280 ;
        RECT 558.630 3.070 559.170 4.280 ;
        RECT 560.010 3.070 560.550 4.280 ;
        RECT 561.390 3.070 561.930 4.280 ;
        RECT 562.770 3.070 563.310 4.280 ;
        RECT 564.150 3.070 564.690 4.280 ;
        RECT 565.530 3.070 566.070 4.280 ;
        RECT 566.910 3.070 567.450 4.280 ;
        RECT 568.290 3.070 568.830 4.280 ;
        RECT 569.670 3.070 570.210 4.280 ;
        RECT 571.050 3.070 571.590 4.280 ;
        RECT 572.430 3.070 572.970 4.280 ;
        RECT 573.810 3.070 574.350 4.280 ;
        RECT 575.190 3.070 575.730 4.280 ;
        RECT 576.570 3.070 577.110 4.280 ;
        RECT 577.950 3.070 578.490 4.280 ;
        RECT 579.330 3.070 579.870 4.280 ;
        RECT 580.710 3.070 581.250 4.280 ;
        RECT 582.090 3.070 582.630 4.280 ;
        RECT 583.470 3.070 584.010 4.280 ;
        RECT 584.850 3.070 585.390 4.280 ;
        RECT 586.230 3.070 586.770 4.280 ;
        RECT 587.610 3.070 588.150 4.280 ;
        RECT 588.990 3.070 589.530 4.280 ;
        RECT 590.370 3.070 590.910 4.280 ;
        RECT 591.750 3.070 592.290 4.280 ;
        RECT 593.130 3.070 593.670 4.280 ;
        RECT 594.510 3.070 595.050 4.280 ;
        RECT 595.890 3.070 596.430 4.280 ;
        RECT 597.270 3.070 597.810 4.280 ;
        RECT 598.650 3.070 599.190 4.280 ;
        RECT 600.030 3.070 600.570 4.280 ;
        RECT 601.410 3.070 601.950 4.280 ;
        RECT 602.790 3.070 603.330 4.280 ;
        RECT 604.170 3.070 604.710 4.280 ;
        RECT 605.550 3.070 606.090 4.280 ;
        RECT 606.930 3.070 607.470 4.280 ;
        RECT 608.310 3.070 608.850 4.280 ;
        RECT 609.690 3.070 610.230 4.280 ;
        RECT 611.070 3.070 611.610 4.280 ;
        RECT 612.450 3.070 612.990 4.280 ;
        RECT 613.830 3.070 614.370 4.280 ;
        RECT 615.210 3.070 615.750 4.280 ;
        RECT 616.590 3.070 617.130 4.280 ;
        RECT 617.970 3.070 618.510 4.280 ;
        RECT 619.350 3.070 619.890 4.280 ;
        RECT 620.730 3.070 621.270 4.280 ;
        RECT 622.110 3.070 622.650 4.280 ;
        RECT 623.490 3.070 624.030 4.280 ;
        RECT 624.870 3.070 625.410 4.280 ;
        RECT 626.250 3.070 626.790 4.280 ;
        RECT 627.630 3.070 628.170 4.280 ;
        RECT 629.010 3.070 629.550 4.280 ;
        RECT 630.390 3.070 630.930 4.280 ;
        RECT 631.770 3.070 632.310 4.280 ;
        RECT 633.150 3.070 633.690 4.280 ;
        RECT 634.530 3.070 635.070 4.280 ;
        RECT 635.910 3.070 636.450 4.280 ;
        RECT 637.290 3.070 637.830 4.280 ;
        RECT 638.670 3.070 639.210 4.280 ;
        RECT 640.050 3.070 640.590 4.280 ;
        RECT 641.430 3.070 641.970 4.280 ;
        RECT 642.810 3.070 643.350 4.280 ;
        RECT 644.190 3.070 644.730 4.280 ;
        RECT 645.570 3.070 646.110 4.280 ;
        RECT 646.950 3.070 647.490 4.280 ;
        RECT 648.330 3.070 648.870 4.280 ;
        RECT 649.710 3.070 650.250 4.280 ;
        RECT 651.090 3.070 651.630 4.280 ;
        RECT 652.470 3.070 653.010 4.280 ;
        RECT 653.850 3.070 654.390 4.280 ;
        RECT 655.230 3.070 655.770 4.280 ;
        RECT 656.610 3.070 657.150 4.280 ;
        RECT 657.990 3.070 658.530 4.280 ;
        RECT 659.370 3.070 659.910 4.280 ;
        RECT 660.750 3.070 661.290 4.280 ;
        RECT 662.130 3.070 662.670 4.280 ;
        RECT 663.510 3.070 664.050 4.280 ;
        RECT 664.890 3.070 665.430 4.280 ;
        RECT 666.270 3.070 666.810 4.280 ;
        RECT 667.650 3.070 668.190 4.280 ;
        RECT 669.030 3.070 669.570 4.280 ;
        RECT 670.410 3.070 670.950 4.280 ;
        RECT 671.790 3.070 672.330 4.280 ;
        RECT 673.170 3.070 673.710 4.280 ;
        RECT 674.550 3.070 675.090 4.280 ;
        RECT 675.930 3.070 676.470 4.280 ;
        RECT 677.310 3.070 677.850 4.280 ;
        RECT 678.690 3.070 679.230 4.280 ;
        RECT 680.070 3.070 680.610 4.280 ;
        RECT 681.450 3.070 681.990 4.280 ;
        RECT 682.830 3.070 683.370 4.280 ;
        RECT 684.210 3.070 684.750 4.280 ;
        RECT 685.590 3.070 686.130 4.280 ;
        RECT 686.970 3.070 687.510 4.280 ;
        RECT 688.350 3.070 688.890 4.280 ;
        RECT 689.730 3.070 690.270 4.280 ;
        RECT 691.110 3.070 691.650 4.280 ;
        RECT 692.490 3.070 693.030 4.280 ;
        RECT 693.870 3.070 694.410 4.280 ;
        RECT 695.250 3.070 695.790 4.280 ;
        RECT 696.630 3.070 697.170 4.280 ;
        RECT 698.010 3.070 698.550 4.280 ;
        RECT 699.390 3.070 699.930 4.280 ;
        RECT 700.770 3.070 701.310 4.280 ;
        RECT 702.150 3.070 702.690 4.280 ;
        RECT 703.530 3.070 704.070 4.280 ;
        RECT 704.910 3.070 705.450 4.280 ;
        RECT 706.290 3.070 706.830 4.280 ;
        RECT 707.670 3.070 708.210 4.280 ;
        RECT 709.050 3.070 709.590 4.280 ;
        RECT 710.430 3.070 710.970 4.280 ;
        RECT 711.810 3.070 712.350 4.280 ;
        RECT 713.190 3.070 713.730 4.280 ;
        RECT 714.570 3.070 715.110 4.280 ;
        RECT 715.950 3.070 716.490 4.280 ;
        RECT 717.330 3.070 717.870 4.280 ;
        RECT 718.710 3.070 719.250 4.280 ;
        RECT 720.090 3.070 720.630 4.280 ;
        RECT 721.470 3.070 722.010 4.280 ;
        RECT 722.850 3.070 723.390 4.280 ;
        RECT 724.230 3.070 724.770 4.280 ;
        RECT 725.610 3.070 726.150 4.280 ;
        RECT 726.990 3.070 727.530 4.280 ;
        RECT 728.370 3.070 728.910 4.280 ;
        RECT 729.750 3.070 730.290 4.280 ;
        RECT 731.130 3.070 731.670 4.280 ;
        RECT 732.510 3.070 733.050 4.280 ;
        RECT 733.890 3.070 734.430 4.280 ;
        RECT 735.270 3.070 735.810 4.280 ;
        RECT 736.650 3.070 737.190 4.280 ;
        RECT 738.030 3.070 738.570 4.280 ;
        RECT 739.410 3.070 739.950 4.280 ;
        RECT 740.790 3.070 741.330 4.280 ;
        RECT 742.170 3.070 742.710 4.280 ;
        RECT 743.550 3.070 744.090 4.280 ;
        RECT 744.930 3.070 745.470 4.280 ;
        RECT 746.310 3.070 746.850 4.280 ;
        RECT 747.690 3.070 748.230 4.280 ;
        RECT 749.070 3.070 749.610 4.280 ;
        RECT 750.450 3.070 750.990 4.280 ;
        RECT 751.830 3.070 752.370 4.280 ;
        RECT 753.210 3.070 753.750 4.280 ;
        RECT 754.590 3.070 755.130 4.280 ;
        RECT 755.970 3.070 756.510 4.280 ;
        RECT 757.350 3.070 757.890 4.280 ;
        RECT 758.730 3.070 759.270 4.280 ;
        RECT 760.110 3.070 760.650 4.280 ;
        RECT 761.490 3.070 762.030 4.280 ;
        RECT 762.870 3.070 763.410 4.280 ;
        RECT 764.250 3.070 764.790 4.280 ;
        RECT 765.630 3.070 766.170 4.280 ;
        RECT 767.010 3.070 767.550 4.280 ;
        RECT 768.390 3.070 768.930 4.280 ;
        RECT 769.770 3.070 770.310 4.280 ;
        RECT 771.150 3.070 771.690 4.280 ;
        RECT 772.530 3.070 773.070 4.280 ;
        RECT 773.910 3.070 774.450 4.280 ;
        RECT 775.290 3.070 775.830 4.280 ;
        RECT 776.670 3.070 777.210 4.280 ;
        RECT 778.050 3.070 778.590 4.280 ;
        RECT 779.430 3.070 779.970 4.280 ;
        RECT 780.810 3.070 781.350 4.280 ;
        RECT 782.190 3.070 782.730 4.280 ;
        RECT 783.570 3.070 784.110 4.280 ;
        RECT 784.950 3.070 785.490 4.280 ;
        RECT 786.330 3.070 786.870 4.280 ;
        RECT 787.710 3.070 788.250 4.280 ;
        RECT 789.090 3.070 789.630 4.280 ;
        RECT 790.470 3.070 891.840 4.280 ;
      LAYER met3 ;
        RECT 21.050 4.935 867.430 587.685 ;
      LAYER met4 ;
        RECT 206.375 10.240 251.040 55.585 ;
        RECT 253.440 10.240 327.840 55.585 ;
        RECT 330.240 10.240 404.640 55.585 ;
        RECT 407.040 10.240 481.440 55.585 ;
        RECT 483.840 10.240 484.545 55.585 ;
        RECT 206.375 4.935 484.545 10.240 ;
  END
END user_proj_example
END LIBRARY


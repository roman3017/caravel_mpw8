// This is the unpowered netlist.
module user_proj_example (user_clock2,
    wb_clk_i,
    wb_rst_i,
    wbs_ack_o,
    wbs_cyc_i,
    wbs_stb_i,
    wbs_we_i,
    io_in,
    io_oeb,
    io_out,
    irq,
    la_data_in,
    la_data_out,
    la_oenb,
    wbs_adr_i,
    wbs_dat_i,
    wbs_dat_o,
    wbs_sel_i);
 input user_clock2;
 input wb_clk_i;
 input wb_rst_i;
 output wbs_ack_o;
 input wbs_cyc_i;
 input wbs_stb_i;
 input wbs_we_i;
 input [37:0] io_in;
 output [37:0] io_oeb;
 output [37:0] io_out;
 output [2:0] irq;
 input [127:0] la_data_in;
 output [127:0] la_data_out;
 input [127:0] la_oenb;
 input [31:0] wbs_adr_i;
 input [31:0] wbs_dat_i;
 output [31:0] wbs_dat_o;
 input [3:0] wbs_sel_i;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire net264;
 wire net265;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net64;
 wire net281;
 wire net266;
 wire net65;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net267;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire clknet_leaf_0_user_clock2;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net66;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net67;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net68;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net113;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net114;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net104;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net105;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net106;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net107;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net108;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net109;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net110;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net111;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net112;
 wire \usb2uart.dn_tx ;
 wire \usb2uart.dp_tx ;
 wire \usb2uart.u_uart.uart_rx_inst.bit_cnt[0] ;
 wire \usb2uart.u_uart.uart_rx_inst.bit_cnt[1] ;
 wire \usb2uart.u_uart.uart_rx_inst.bit_cnt[2] ;
 wire \usb2uart.u_uart.uart_rx_inst.bit_cnt[3] ;
 wire \usb2uart.u_uart.uart_rx_inst.data_reg[0] ;
 wire \usb2uart.u_uart.uart_rx_inst.data_reg[1] ;
 wire \usb2uart.u_uart.uart_rx_inst.data_reg[2] ;
 wire \usb2uart.u_uart.uart_rx_inst.data_reg[3] ;
 wire \usb2uart.u_uart.uart_rx_inst.data_reg[4] ;
 wire \usb2uart.u_uart.uart_rx_inst.data_reg[5] ;
 wire \usb2uart.u_uart.uart_rx_inst.data_reg[6] ;
 wire \usb2uart.u_uart.uart_rx_inst.data_reg[7] ;
 wire \usb2uart.u_uart.uart_rx_inst.m_axis_tdata_reg[0] ;
 wire \usb2uart.u_uart.uart_rx_inst.m_axis_tdata_reg[1] ;
 wire \usb2uart.u_uart.uart_rx_inst.m_axis_tdata_reg[2] ;
 wire \usb2uart.u_uart.uart_rx_inst.m_axis_tdata_reg[3] ;
 wire \usb2uart.u_uart.uart_rx_inst.m_axis_tdata_reg[4] ;
 wire \usb2uart.u_uart.uart_rx_inst.m_axis_tdata_reg[5] ;
 wire \usb2uart.u_uart.uart_rx_inst.m_axis_tdata_reg[6] ;
 wire \usb2uart.u_uart.uart_rx_inst.m_axis_tdata_reg[7] ;
 wire \usb2uart.u_uart.uart_rx_inst.m_axis_tvalid_reg ;
 wire \usb2uart.u_uart.uart_rx_inst.prescale_reg[0] ;
 wire \usb2uart.u_uart.uart_rx_inst.prescale_reg[10] ;
 wire \usb2uart.u_uart.uart_rx_inst.prescale_reg[11] ;
 wire \usb2uart.u_uart.uart_rx_inst.prescale_reg[12] ;
 wire \usb2uart.u_uart.uart_rx_inst.prescale_reg[13] ;
 wire \usb2uart.u_uart.uart_rx_inst.prescale_reg[14] ;
 wire \usb2uart.u_uart.uart_rx_inst.prescale_reg[15] ;
 wire \usb2uart.u_uart.uart_rx_inst.prescale_reg[16] ;
 wire \usb2uart.u_uart.uart_rx_inst.prescale_reg[17] ;
 wire \usb2uart.u_uart.uart_rx_inst.prescale_reg[18] ;
 wire \usb2uart.u_uart.uart_rx_inst.prescale_reg[1] ;
 wire \usb2uart.u_uart.uart_rx_inst.prescale_reg[2] ;
 wire \usb2uart.u_uart.uart_rx_inst.prescale_reg[3] ;
 wire \usb2uart.u_uart.uart_rx_inst.prescale_reg[4] ;
 wire \usb2uart.u_uart.uart_rx_inst.prescale_reg[5] ;
 wire \usb2uart.u_uart.uart_rx_inst.prescale_reg[6] ;
 wire \usb2uart.u_uart.uart_rx_inst.prescale_reg[7] ;
 wire \usb2uart.u_uart.uart_rx_inst.prescale_reg[8] ;
 wire \usb2uart.u_uart.uart_rx_inst.prescale_reg[9] ;
 wire \usb2uart.u_uart.uart_rx_inst.rxd_reg ;
 wire \usb2uart.u_uart.uart_tx_inst.bit_cnt[0] ;
 wire \usb2uart.u_uart.uart_tx_inst.bit_cnt[1] ;
 wire \usb2uart.u_uart.uart_tx_inst.bit_cnt[2] ;
 wire \usb2uart.u_uart.uart_tx_inst.bit_cnt[3] ;
 wire \usb2uart.u_uart.uart_tx_inst.data_reg[0] ;
 wire \usb2uart.u_uart.uart_tx_inst.data_reg[1] ;
 wire \usb2uart.u_uart.uart_tx_inst.data_reg[2] ;
 wire \usb2uart.u_uart.uart_tx_inst.data_reg[3] ;
 wire \usb2uart.u_uart.uart_tx_inst.data_reg[4] ;
 wire \usb2uart.u_uart.uart_tx_inst.data_reg[5] ;
 wire \usb2uart.u_uart.uart_tx_inst.data_reg[6] ;
 wire \usb2uart.u_uart.uart_tx_inst.data_reg[7] ;
 wire \usb2uart.u_uart.uart_tx_inst.data_reg[8] ;
 wire \usb2uart.u_uart.uart_tx_inst.prescale_reg[0] ;
 wire \usb2uart.u_uart.uart_tx_inst.prescale_reg[10] ;
 wire \usb2uart.u_uart.uart_tx_inst.prescale_reg[11] ;
 wire \usb2uart.u_uart.uart_tx_inst.prescale_reg[12] ;
 wire \usb2uart.u_uart.uart_tx_inst.prescale_reg[13] ;
 wire \usb2uart.u_uart.uart_tx_inst.prescale_reg[14] ;
 wire \usb2uart.u_uart.uart_tx_inst.prescale_reg[15] ;
 wire \usb2uart.u_uart.uart_tx_inst.prescale_reg[16] ;
 wire \usb2uart.u_uart.uart_tx_inst.prescale_reg[17] ;
 wire \usb2uart.u_uart.uart_tx_inst.prescale_reg[18] ;
 wire \usb2uart.u_uart.uart_tx_inst.prescale_reg[1] ;
 wire \usb2uart.u_uart.uart_tx_inst.prescale_reg[2] ;
 wire \usb2uart.u_uart.uart_tx_inst.prescale_reg[3] ;
 wire \usb2uart.u_uart.uart_tx_inst.prescale_reg[4] ;
 wire \usb2uart.u_uart.uart_tx_inst.prescale_reg[5] ;
 wire \usb2uart.u_uart.uart_tx_inst.prescale_reg[6] ;
 wire \usb2uart.u_uart.uart_tx_inst.prescale_reg[7] ;
 wire \usb2uart.u_uart.uart_tx_inst.prescale_reg[8] ;
 wire \usb2uart.u_uart.uart_tx_inst.prescale_reg[9] ;
 wire \usb2uart.u_uart.uart_tx_inst.s_axis_tready_reg ;
 wire \usb2uart.u_usb_cdc.addr[0] ;
 wire \usb2uart.u_usb_cdc.addr[1] ;
 wire \usb2uart.u_usb_cdc.addr[2] ;
 wire \usb2uart.u_usb_cdc.addr[3] ;
 wire \usb2uart.u_usb_cdc.addr[4] ;
 wire \usb2uart.u_usb_cdc.addr[5] ;
 wire \usb2uart.u_usb_cdc.addr[6] ;
 wire \usb2uart.u_usb_cdc.bulk_in_req ;
 wire \usb2uart.u_usb_cdc.bulk_in_valid ;
 wire \usb2uart.u_usb_cdc.bulk_out_nak ;
 wire \usb2uart.u_usb_cdc.ctrl_in_req ;
 wire \usb2uart.u_usb_cdc.ctrl_stall ;
 wire \usb2uart.u_usb_cdc.endp[0] ;
 wire \usb2uart.u_usb_cdc.endp[1] ;
 wire \usb2uart.u_usb_cdc.endp[2] ;
 wire \usb2uart.u_usb_cdc.endp[3] ;
 wire \usb2uart.u_usb_cdc.in_data_ack ;
 wire \usb2uart.u_usb_cdc.out_data[0] ;
 wire \usb2uart.u_usb_cdc.out_data[1] ;
 wire \usb2uart.u_usb_cdc.out_data[2] ;
 wire \usb2uart.u_usb_cdc.out_data[3] ;
 wire \usb2uart.u_usb_cdc.out_data[4] ;
 wire \usb2uart.u_usb_cdc.out_data[5] ;
 wire \usb2uart.u_usb_cdc.out_data[6] ;
 wire \usb2uart.u_usb_cdc.out_data[7] ;
 wire \usb2uart.u_usb_cdc.out_err ;
 wire \usb2uart.u_usb_cdc.rstn ;
 wire \usb2uart.u_usb_cdc.rstn_sq[1] ;
 wire \usb2uart.u_usb_cdc.u_bulk_endp.rstn ;
 wire \usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.delay_in_cnt_q[0] ;
 wire \usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.delay_in_cnt_q[1] ;
 wire \usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[0] ;
 wire \usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[10] ;
 wire \usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[11] ;
 wire \usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[12] ;
 wire \usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[13] ;
 wire \usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[14] ;
 wire \usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[15] ;
 wire \usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[16] ;
 wire \usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[17] ;
 wire \usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[18] ;
 wire \usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[19] ;
 wire \usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[1] ;
 wire \usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[20] ;
 wire \usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[21] ;
 wire \usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[22] ;
 wire \usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[23] ;
 wire \usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[24] ;
 wire \usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[25] ;
 wire \usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[26] ;
 wire \usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[27] ;
 wire \usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[28] ;
 wire \usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[29] ;
 wire \usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[2] ;
 wire \usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[30] ;
 wire \usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[31] ;
 wire \usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[32] ;
 wire \usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[33] ;
 wire \usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[34] ;
 wire \usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[35] ;
 wire \usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[36] ;
 wire \usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[37] ;
 wire \usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[38] ;
 wire \usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[39] ;
 wire \usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[3] ;
 wire \usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[40] ;
 wire \usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[41] ;
 wire \usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[42] ;
 wire \usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[43] ;
 wire \usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[44] ;
 wire \usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[45] ;
 wire \usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[46] ;
 wire \usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[47] ;
 wire \usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[48] ;
 wire \usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[49] ;
 wire \usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[4] ;
 wire \usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[50] ;
 wire \usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[51] ;
 wire \usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[52] ;
 wire \usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[53] ;
 wire \usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[54] ;
 wire \usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[55] ;
 wire \usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[56] ;
 wire \usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[57] ;
 wire \usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[58] ;
 wire \usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[59] ;
 wire \usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[5] ;
 wire \usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[60] ;
 wire \usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[61] ;
 wire \usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[62] ;
 wire \usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[63] ;
 wire \usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[64] ;
 wire \usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[65] ;
 wire \usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[66] ;
 wire \usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[67] ;
 wire \usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[68] ;
 wire \usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[69] ;
 wire \usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[6] ;
 wire \usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[70] ;
 wire \usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[71] ;
 wire \usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[7] ;
 wire \usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[8] ;
 wire \usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[9] ;
 wire \usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_first_q[0] ;
 wire \usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_first_q[1] ;
 wire \usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_first_q[2] ;
 wire \usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_first_q[3] ;
 wire \usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_first_qq[0] ;
 wire \usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_first_qq[1] ;
 wire \usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_first_qq[2] ;
 wire \usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_first_qq[3] ;
 wire \usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_last_q[0] ;
 wire \usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_last_q[1] ;
 wire \usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_last_q[2] ;
 wire \usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_last_q[3] ;
 wire \usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_req_q ;
 wire \usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_state_q ;
 wire \usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.delay_out_cnt_q[0] ;
 wire \usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.delay_out_cnt_q[1] ;
 wire \usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[0] ;
 wire \usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[10] ;
 wire \usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[11] ;
 wire \usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[12] ;
 wire \usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[13] ;
 wire \usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[14] ;
 wire \usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[15] ;
 wire \usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[16] ;
 wire \usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[17] ;
 wire \usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[18] ;
 wire \usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[19] ;
 wire \usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[1] ;
 wire \usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[20] ;
 wire \usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[21] ;
 wire \usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[22] ;
 wire \usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[23] ;
 wire \usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[24] ;
 wire \usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[25] ;
 wire \usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[26] ;
 wire \usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[27] ;
 wire \usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[28] ;
 wire \usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[29] ;
 wire \usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[2] ;
 wire \usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[30] ;
 wire \usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[31] ;
 wire \usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[32] ;
 wire \usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[33] ;
 wire \usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[34] ;
 wire \usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[35] ;
 wire \usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[36] ;
 wire \usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[37] ;
 wire \usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[38] ;
 wire \usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[39] ;
 wire \usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[3] ;
 wire \usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[40] ;
 wire \usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[41] ;
 wire \usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[42] ;
 wire \usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[43] ;
 wire \usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[44] ;
 wire \usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[45] ;
 wire \usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[46] ;
 wire \usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[47] ;
 wire \usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[48] ;
 wire \usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[49] ;
 wire \usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[4] ;
 wire \usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[50] ;
 wire \usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[51] ;
 wire \usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[52] ;
 wire \usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[53] ;
 wire \usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[54] ;
 wire \usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[55] ;
 wire \usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[56] ;
 wire \usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[57] ;
 wire \usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[58] ;
 wire \usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[59] ;
 wire \usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[5] ;
 wire \usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[60] ;
 wire \usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[61] ;
 wire \usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[62] ;
 wire \usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[63] ;
 wire \usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[64] ;
 wire \usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[65] ;
 wire \usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[66] ;
 wire \usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[67] ;
 wire \usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[68] ;
 wire \usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[69] ;
 wire \usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[6] ;
 wire \usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[70] ;
 wire \usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[71] ;
 wire \usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[7] ;
 wire \usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[8] ;
 wire \usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[9] ;
 wire \usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_first_q[0] ;
 wire \usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_first_q[1] ;
 wire \usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_first_q[2] ;
 wire \usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_first_q[3] ;
 wire \usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_full_o ;
 wire \usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_last_q[0] ;
 wire \usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_last_q[1] ;
 wire \usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_last_q[2] ;
 wire \usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_last_q[3] ;
 wire \usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_last_qq[0] ;
 wire \usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_last_qq[1] ;
 wire \usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_last_qq[2] ;
 wire \usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_last_qq[3] ;
 wire \usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_state_q[1] ;
 wire \usb2uart.u_usb_cdc.u_ctrl_endp.addr_q[0] ;
 wire \usb2uart.u_usb_cdc.u_ctrl_endp.addr_q[1] ;
 wire \usb2uart.u_usb_cdc.u_ctrl_endp.addr_q[2] ;
 wire \usb2uart.u_usb_cdc.u_ctrl_endp.addr_q[3] ;
 wire \usb2uart.u_usb_cdc.u_ctrl_endp.addr_q[4] ;
 wire \usb2uart.u_usb_cdc.u_ctrl_endp.addr_q[5] ;
 wire \usb2uart.u_usb_cdc.u_ctrl_endp.addr_q[6] ;
 wire \usb2uart.u_usb_cdc.u_ctrl_endp.byte_cnt_q[0] ;
 wire \usb2uart.u_usb_cdc.u_ctrl_endp.byte_cnt_q[1] ;
 wire \usb2uart.u_usb_cdc.u_ctrl_endp.byte_cnt_q[2] ;
 wire \usb2uart.u_usb_cdc.u_ctrl_endp.byte_cnt_q[3] ;
 wire \usb2uart.u_usb_cdc.u_ctrl_endp.byte_cnt_q[4] ;
 wire \usb2uart.u_usb_cdc.u_ctrl_endp.byte_cnt_q[5] ;
 wire \usb2uart.u_usb_cdc.u_ctrl_endp.byte_cnt_q[6] ;
 wire \usb2uart.u_usb_cdc.u_ctrl_endp.class_q ;
 wire \usb2uart.u_usb_cdc.u_ctrl_endp.dev_state_q[0] ;
 wire \usb2uart.u_usb_cdc.u_ctrl_endp.dev_state_q[1] ;
 wire \usb2uart.u_usb_cdc.u_ctrl_endp.dev_state_qq[0] ;
 wire \usb2uart.u_usb_cdc.u_ctrl_endp.dev_state_qq[1] ;
 wire \usb2uart.u_usb_cdc.u_ctrl_endp.in_dir_q ;
 wire \usb2uart.u_usb_cdc.u_ctrl_endp.in_endp_q ;
 wire \usb2uart.u_usb_cdc.u_ctrl_endp.in_req_q ;
 wire \usb2uart.u_usb_cdc.u_ctrl_endp.max_length_q[0] ;
 wire \usb2uart.u_usb_cdc.u_ctrl_endp.max_length_q[1] ;
 wire \usb2uart.u_usb_cdc.u_ctrl_endp.max_length_q[2] ;
 wire \usb2uart.u_usb_cdc.u_ctrl_endp.max_length_q[3] ;
 wire \usb2uart.u_usb_cdc.u_ctrl_endp.max_length_q[4] ;
 wire \usb2uart.u_usb_cdc.u_ctrl_endp.max_length_q[5] ;
 wire \usb2uart.u_usb_cdc.u_ctrl_endp.max_length_q[6] ;
 wire \usb2uart.u_usb_cdc.u_ctrl_endp.rec_q[0] ;
 wire \usb2uart.u_usb_cdc.u_ctrl_endp.rec_q[1] ;
 wire \usb2uart.u_usb_cdc.u_ctrl_endp.req_q[0] ;
 wire \usb2uart.u_usb_cdc.u_ctrl_endp.req_q[10] ;
 wire \usb2uart.u_usb_cdc.u_ctrl_endp.req_q[11] ;
 wire \usb2uart.u_usb_cdc.u_ctrl_endp.req_q[1] ;
 wire \usb2uart.u_usb_cdc.u_ctrl_endp.req_q[2] ;
 wire \usb2uart.u_usb_cdc.u_ctrl_endp.req_q[3] ;
 wire \usb2uart.u_usb_cdc.u_ctrl_endp.req_q[4] ;
 wire \usb2uart.u_usb_cdc.u_ctrl_endp.req_q[5] ;
 wire \usb2uart.u_usb_cdc.u_ctrl_endp.req_q[6] ;
 wire \usb2uart.u_usb_cdc.u_ctrl_endp.req_q[7] ;
 wire \usb2uart.u_usb_cdc.u_ctrl_endp.req_q[8] ;
 wire \usb2uart.u_usb_cdc.u_ctrl_endp.req_q[9] ;
 wire \usb2uart.u_usb_cdc.u_ctrl_endp.state_q[0] ;
 wire \usb2uart.u_usb_cdc.u_ctrl_endp.state_q[1] ;
 wire \usb2uart.u_usb_cdc.u_ctrl_endp.state_q[3] ;
 wire \usb2uart.u_usb_cdc.u_ctrl_endp.usb_reset_q ;
 wire \usb2uart.u_usb_cdc.u_sie.addr_q[0] ;
 wire \usb2uart.u_usb_cdc.u_sie.addr_q[1] ;
 wire \usb2uart.u_usb_cdc.u_sie.addr_q[2] ;
 wire \usb2uart.u_usb_cdc.u_sie.addr_q[3] ;
 wire \usb2uart.u_usb_cdc.u_sie.addr_q[4] ;
 wire \usb2uart.u_usb_cdc.u_sie.addr_q[5] ;
 wire \usb2uart.u_usb_cdc.u_sie.addr_q[6] ;
 wire \usb2uart.u_usb_cdc.u_sie.crc16_q[0] ;
 wire \usb2uart.u_usb_cdc.u_sie.crc16_q[10] ;
 wire \usb2uart.u_usb_cdc.u_sie.crc16_q[11] ;
 wire \usb2uart.u_usb_cdc.u_sie.crc16_q[12] ;
 wire \usb2uart.u_usb_cdc.u_sie.crc16_q[13] ;
 wire \usb2uart.u_usb_cdc.u_sie.crc16_q[14] ;
 wire \usb2uart.u_usb_cdc.u_sie.crc16_q[15] ;
 wire \usb2uart.u_usb_cdc.u_sie.crc16_q[1] ;
 wire \usb2uart.u_usb_cdc.u_sie.crc16_q[2] ;
 wire \usb2uart.u_usb_cdc.u_sie.crc16_q[3] ;
 wire \usb2uart.u_usb_cdc.u_sie.crc16_q[4] ;
 wire \usb2uart.u_usb_cdc.u_sie.crc16_q[5] ;
 wire \usb2uart.u_usb_cdc.u_sie.crc16_q[6] ;
 wire \usb2uart.u_usb_cdc.u_sie.crc16_q[7] ;
 wire \usb2uart.u_usb_cdc.u_sie.crc16_q[8] ;
 wire \usb2uart.u_usb_cdc.u_sie.crc16_q[9] ;
 wire \usb2uart.u_usb_cdc.u_sie.data_q[0] ;
 wire \usb2uart.u_usb_cdc.u_sie.data_q[1] ;
 wire \usb2uart.u_usb_cdc.u_sie.data_q[2] ;
 wire \usb2uart.u_usb_cdc.u_sie.data_q[3] ;
 wire \usb2uart.u_usb_cdc.u_sie.data_q[4] ;
 wire \usb2uart.u_usb_cdc.u_sie.data_q[5] ;
 wire \usb2uart.u_usb_cdc.u_sie.data_q[6] ;
 wire \usb2uart.u_usb_cdc.u_sie.data_q[7] ;
 wire \usb2uart.u_usb_cdc.u_sie.datain_toggle_q[0] ;
 wire \usb2uart.u_usb_cdc.u_sie.datain_toggle_q[1] ;
 wire \usb2uart.u_usb_cdc.u_sie.dataout_toggle_q[0] ;
 wire \usb2uart.u_usb_cdc.u_sie.dataout_toggle_q[1] ;
 wire \usb2uart.u_usb_cdc.u_sie.delay_cnt_q[0] ;
 wire \usb2uart.u_usb_cdc.u_sie.delay_cnt_q[1] ;
 wire \usb2uart.u_usb_cdc.u_sie.delay_cnt_q[2] ;
 wire \usb2uart.u_usb_cdc.u_sie.delay_cnt_q[3] ;
 wire \usb2uart.u_usb_cdc.u_sie.delay_cnt_q[4] ;
 wire \usb2uart.u_usb_cdc.u_sie.in_byte_q[0] ;
 wire \usb2uart.u_usb_cdc.u_sie.in_byte_q[1] ;
 wire \usb2uart.u_usb_cdc.u_sie.in_byte_q[2] ;
 wire \usb2uart.u_usb_cdc.u_sie.in_byte_q[3] ;
 wire \usb2uart.u_usb_cdc.u_sie.out_eop_q ;
 wire \usb2uart.u_usb_cdc.u_sie.phy_state_q[0] ;
 wire \usb2uart.u_usb_cdc.u_sie.phy_state_q[10] ;
 wire \usb2uart.u_usb_cdc.u_sie.phy_state_q[11] ;
 wire \usb2uart.u_usb_cdc.u_sie.phy_state_q[1] ;
 wire \usb2uart.u_usb_cdc.u_sie.phy_state_q[2] ;
 wire \usb2uart.u_usb_cdc.u_sie.phy_state_q[3] ;
 wire \usb2uart.u_usb_cdc.u_sie.phy_state_q[4] ;
 wire \usb2uart.u_usb_cdc.u_sie.phy_state_q[5] ;
 wire \usb2uart.u_usb_cdc.u_sie.phy_state_q[6] ;
 wire \usb2uart.u_usb_cdc.u_sie.phy_state_q[7] ;
 wire \usb2uart.u_usb_cdc.u_sie.phy_state_q[8] ;
 wire \usb2uart.u_usb_cdc.u_sie.phy_state_q[9] ;
 wire \usb2uart.u_usb_cdc.u_sie.pid_q[0] ;
 wire \usb2uart.u_usb_cdc.u_sie.pid_q[1] ;
 wire \usb2uart.u_usb_cdc.u_sie.pid_q[2] ;
 wire \usb2uart.u_usb_cdc.u_sie.pid_q[3] ;
 wire \usb2uart.u_usb_cdc.u_sie.rx_data[0] ;
 wire \usb2uart.u_usb_cdc.u_sie.rx_data[1] ;
 wire \usb2uart.u_usb_cdc.u_sie.rx_data[2] ;
 wire \usb2uart.u_usb_cdc.u_sie.rx_data[3] ;
 wire \usb2uart.u_usb_cdc.u_sie.rx_data[4] ;
 wire \usb2uart.u_usb_cdc.u_sie.rx_data[5] ;
 wire \usb2uart.u_usb_cdc.u_sie.rx_data[6] ;
 wire \usb2uart.u_usb_cdc.u_sie.rx_data[7] ;
 wire \usb2uart.u_usb_cdc.u_sie.rx_err ;
 wire \usb2uart.u_usb_cdc.u_sie.u_phy_rx.clk_cnt_q[0] ;
 wire \usb2uart.u_usb_cdc.u_sie.u_phy_rx.clk_cnt_q[1] ;
 wire \usb2uart.u_usb_cdc.u_sie.u_phy_rx.cnt_q[0] ;
 wire \usb2uart.u_usb_cdc.u_sie.u_phy_rx.cnt_q[10] ;
 wire \usb2uart.u_usb_cdc.u_sie.u_phy_rx.cnt_q[11] ;
 wire \usb2uart.u_usb_cdc.u_sie.u_phy_rx.cnt_q[12] ;
 wire \usb2uart.u_usb_cdc.u_sie.u_phy_rx.cnt_q[13] ;
 wire \usb2uart.u_usb_cdc.u_sie.u_phy_rx.cnt_q[14] ;
 wire \usb2uart.u_usb_cdc.u_sie.u_phy_rx.cnt_q[15] ;
 wire \usb2uart.u_usb_cdc.u_sie.u_phy_rx.cnt_q[16] ;
 wire \usb2uart.u_usb_cdc.u_sie.u_phy_rx.cnt_q[17] ;
 wire \usb2uart.u_usb_cdc.u_sie.u_phy_rx.cnt_q[1] ;
 wire \usb2uart.u_usb_cdc.u_sie.u_phy_rx.cnt_q[2] ;
 wire \usb2uart.u_usb_cdc.u_sie.u_phy_rx.cnt_q[3] ;
 wire \usb2uart.u_usb_cdc.u_sie.u_phy_rx.cnt_q[4] ;
 wire \usb2uart.u_usb_cdc.u_sie.u_phy_rx.cnt_q[5] ;
 wire \usb2uart.u_usb_cdc.u_sie.u_phy_rx.cnt_q[6] ;
 wire \usb2uart.u_usb_cdc.u_sie.u_phy_rx.cnt_q[7] ;
 wire \usb2uart.u_usb_cdc.u_sie.u_phy_rx.cnt_q[8] ;
 wire \usb2uart.u_usb_cdc.u_sie.u_phy_rx.cnt_q[9] ;
 wire \usb2uart.u_usb_cdc.u_sie.u_phy_rx.data_q[0] ;
 wire \usb2uart.u_usb_cdc.u_sie.u_phy_rx.dn_q[0] ;
 wire \usb2uart.u_usb_cdc.u_sie.u_phy_rx.dn_q[1] ;
 wire \usb2uart.u_usb_cdc.u_sie.u_phy_rx.dn_q[2] ;
 wire \usb2uart.u_usb_cdc.u_sie.u_phy_rx.dp_q[0] ;
 wire \usb2uart.u_usb_cdc.u_sie.u_phy_rx.dp_q[1] ;
 wire \usb2uart.u_usb_cdc.u_sie.u_phy_rx.dp_q[2] ;
 wire \usb2uart.u_usb_cdc.u_sie.u_phy_rx.nrzi_q[0] ;
 wire \usb2uart.u_usb_cdc.u_sie.u_phy_rx.nrzi_q[1] ;
 wire \usb2uart.u_usb_cdc.u_sie.u_phy_rx.nrzi_q[2] ;
 wire \usb2uart.u_usb_cdc.u_sie.u_phy_rx.nrzi_q[3] ;
 wire \usb2uart.u_usb_cdc.u_sie.u_phy_rx.rx_en_q ;
 wire \usb2uart.u_usb_cdc.u_sie.u_phy_rx.rx_state_q[0] ;
 wire \usb2uart.u_usb_cdc.u_sie.u_phy_rx.rx_state_q[2] ;
 wire \usb2uart.u_usb_cdc.u_sie.u_phy_rx.rx_state_q[3] ;
 wire \usb2uart.u_usb_cdc.u_sie.u_phy_rx.rx_state_q[4] ;
 wire \usb2uart.u_usb_cdc.u_sie.u_phy_rx.rx_valid_fd ;
 wire \usb2uart.u_usb_cdc.u_sie.u_phy_rx.rx_valid_fq ;
 wire \usb2uart.u_usb_cdc.u_sie.u_phy_rx.stuffing_cnt_q[0] ;
 wire \usb2uart.u_usb_cdc.u_sie.u_phy_rx.stuffing_cnt_q[1] ;
 wire \usb2uart.u_usb_cdc.u_sie.u_phy_rx.stuffing_cnt_q[2] ;
 wire \usb2uart.u_usb_cdc.u_sie.u_phy_tx.bit_cnt_q[0] ;
 wire \usb2uart.u_usb_cdc.u_sie.u_phy_tx.bit_cnt_q[1] ;
 wire \usb2uart.u_usb_cdc.u_sie.u_phy_tx.bit_cnt_q[2] ;
 wire \usb2uart.u_usb_cdc.u_sie.u_phy_tx.clk_cnt_q[0] ;
 wire \usb2uart.u_usb_cdc.u_sie.u_phy_tx.clk_cnt_q[1] ;
 wire \usb2uart.u_usb_cdc.u_sie.u_phy_tx.data_q[0] ;
 wire \usb2uart.u_usb_cdc.u_sie.u_phy_tx.data_q[1] ;
 wire \usb2uart.u_usb_cdc.u_sie.u_phy_tx.data_q[2] ;
 wire \usb2uart.u_usb_cdc.u_sie.u_phy_tx.data_q[3] ;
 wire \usb2uart.u_usb_cdc.u_sie.u_phy_tx.data_q[4] ;
 wire \usb2uart.u_usb_cdc.u_sie.u_phy_tx.data_q[5] ;
 wire \usb2uart.u_usb_cdc.u_sie.u_phy_tx.data_q[6] ;
 wire \usb2uart.u_usb_cdc.u_sie.u_phy_tx.data_q[7] ;
 wire \usb2uart.u_usb_cdc.u_sie.u_phy_tx.nrzi_q ;
 wire \usb2uart.u_usb_cdc.u_sie.u_phy_tx.stuffing_cnt_q[0] ;
 wire \usb2uart.u_usb_cdc.u_sie.u_phy_tx.stuffing_cnt_q[1] ;
 wire \usb2uart.u_usb_cdc.u_sie.u_phy_tx.stuffing_cnt_q[2] ;
 wire \usb2uart.u_usb_cdc.u_sie.u_phy_tx.tx_state_q[1] ;
 wire \usb2uart.u_usb_cdc.u_sie.u_phy_tx.tx_state_q[2] ;
 wire \usb2uart.u_usb_cdc.u_sie.u_phy_tx.tx_state_q[3] ;
 wire \usb2uart.u_usb_cdc.u_sie.u_phy_tx.tx_valid_q ;
 wire net231;
 wire net232;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net233;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net234;
 wire net262;
 wire net263;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire clknet_leaf_1_user_clock2;
 wire clknet_leaf_2_user_clock2;
 wire clknet_leaf_3_user_clock2;
 wire clknet_leaf_4_user_clock2;
 wire clknet_leaf_5_user_clock2;
 wire clknet_leaf_6_user_clock2;
 wire clknet_leaf_8_user_clock2;
 wire clknet_leaf_9_user_clock2;
 wire clknet_leaf_10_user_clock2;
 wire clknet_leaf_11_user_clock2;
 wire clknet_leaf_12_user_clock2;
 wire clknet_leaf_13_user_clock2;
 wire clknet_leaf_14_user_clock2;
 wire clknet_leaf_15_user_clock2;
 wire clknet_leaf_16_user_clock2;
 wire clknet_leaf_17_user_clock2;
 wire clknet_leaf_18_user_clock2;
 wire clknet_leaf_19_user_clock2;
 wire clknet_leaf_20_user_clock2;
 wire clknet_leaf_21_user_clock2;
 wire clknet_leaf_22_user_clock2;
 wire clknet_leaf_23_user_clock2;
 wire clknet_leaf_24_user_clock2;
 wire clknet_leaf_25_user_clock2;
 wire clknet_leaf_26_user_clock2;
 wire clknet_leaf_27_user_clock2;
 wire clknet_leaf_28_user_clock2;
 wire clknet_leaf_29_user_clock2;
 wire clknet_leaf_30_user_clock2;
 wire clknet_leaf_31_user_clock2;
 wire clknet_leaf_32_user_clock2;
 wire clknet_leaf_33_user_clock2;
 wire clknet_leaf_34_user_clock2;
 wire clknet_leaf_35_user_clock2;
 wire clknet_leaf_36_user_clock2;
 wire clknet_leaf_37_user_clock2;
 wire clknet_0_user_clock2;
 wire clknet_2_0__leaf_user_clock2;
 wire clknet_2_1__leaf_user_clock2;
 wire clknet_2_2__leaf_user_clock2;
 wire clknet_2_3__leaf_user_clock2;
 wire clknet_opt_1_0_user_clock2;
 wire net298;
 wire net299;
 wire net300;
 wire net301;

 sky130_fd_sc_hd__clkbuf_1 _2088_ (.A(net6),
    .X(_2001_));
 sky130_fd_sc_hd__clkbuf_1 _2089_ (.A(_2001_),
    .X(_2085_));
 sky130_fd_sc_hd__inv_2 _2090_ (.A(\usb2uart.u_usb_cdc.u_ctrl_endp.class_q ),
    .Y(_2002_));
 sky130_fd_sc_hd__inv_2 _2091_ (.A(\usb2uart.u_usb_cdc.u_sie.rx_err ),
    .Y(_2003_));
 sky130_fd_sc_hd__xor2_4 _2092_ (.A(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.rx_valid_fq ),
    .B(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.rx_valid_fd ),
    .X(_2004_));
 sky130_fd_sc_hd__and3_1 _2093_ (.A(_2003_),
    .B(\usb2uart.u_usb_cdc.u_sie.phy_state_q[8] ),
    .C(_2004_),
    .X(_2005_));
 sky130_fd_sc_hd__buf_2 _2094_ (.A(_2005_),
    .X(_2006_));
 sky130_fd_sc_hd__nor3_2 _2095_ (.A(\usb2uart.u_usb_cdc.endp[1] ),
    .B(\usb2uart.u_usb_cdc.endp[3] ),
    .C(\usb2uart.u_usb_cdc.endp[2] ),
    .Y(_2007_));
 sky130_fd_sc_hd__and2b_1 _2096_ (.A_N(\usb2uart.u_usb_cdc.endp[0] ),
    .B(_2007_),
    .X(_2008_));
 sky130_fd_sc_hd__buf_2 _2097_ (.A(_2008_),
    .X(_2009_));
 sky130_fd_sc_hd__and2b_1 _2098_ (.A_N(\usb2uart.u_usb_cdc.u_ctrl_endp.in_dir_q ),
    .B(\usb2uart.u_usb_cdc.u_ctrl_endp.state_q[3] ),
    .X(_2010_));
 sky130_fd_sc_hd__inv_2 _2099_ (.A(_2010_),
    .Y(_2011_));
 sky130_fd_sc_hd__clkinv_2 _2100_ (.A(\usb2uart.u_usb_cdc.u_ctrl_endp.state_q[1] ),
    .Y(_2012_));
 sky130_fd_sc_hd__or4_1 _2101_ (.A(\usb2uart.u_usb_cdc.u_ctrl_endp.max_length_q[0] ),
    .B(\usb2uart.u_usb_cdc.u_ctrl_endp.max_length_q[1] ),
    .C(\usb2uart.u_usb_cdc.u_ctrl_endp.max_length_q[2] ),
    .D(\usb2uart.u_usb_cdc.u_ctrl_endp.max_length_q[3] ),
    .X(_2013_));
 sky130_fd_sc_hd__or4_1 _2102_ (.A(\usb2uart.u_usb_cdc.u_ctrl_endp.max_length_q[4] ),
    .B(\usb2uart.u_usb_cdc.u_ctrl_endp.max_length_q[5] ),
    .C(\usb2uart.u_usb_cdc.u_ctrl_endp.max_length_q[6] ),
    .D(\usb2uart.u_usb_cdc.u_ctrl_endp.in_dir_q ),
    .X(_2014_));
 sky130_fd_sc_hd__or4b_2 _2103_ (.A(\usb2uart.u_usb_cdc.u_ctrl_endp.byte_cnt_q[2] ),
    .B(\usb2uart.u_usb_cdc.u_ctrl_endp.byte_cnt_q[4] ),
    .C(\usb2uart.u_usb_cdc.u_ctrl_endp.byte_cnt_q[5] ),
    .D_N(\usb2uart.u_usb_cdc.u_ctrl_endp.byte_cnt_q[3] ),
    .X(_2015_));
 sky130_fd_sc_hd__or4_1 _2104_ (.A(\usb2uart.u_usb_cdc.u_ctrl_endp.byte_cnt_q[0] ),
    .B(\usb2uart.u_usb_cdc.u_ctrl_endp.byte_cnt_q[1] ),
    .C(\usb2uart.u_usb_cdc.u_ctrl_endp.byte_cnt_q[6] ),
    .D(\usb2uart.u_usb_cdc.u_ctrl_endp.req_q[10] ),
    .X(_2016_));
 sky130_fd_sc_hd__or4_4 _2105_ (.A(_2013_),
    .B(_2014_),
    .C(_2015_),
    .D(_2016_),
    .X(_2017_));
 sky130_fd_sc_hd__or3_1 _2106_ (.A(_2012_),
    .B(_2005_),
    .C(_2017_),
    .X(_2018_));
 sky130_fd_sc_hd__and4b_1 _2107_ (.A_N(\usb2uart.u_usb_cdc.u_sie.pid_q[1] ),
    .B(\usb2uart.u_usb_cdc.u_sie.pid_q[3] ),
    .C(\usb2uart.u_usb_cdc.u_sie.pid_q[2] ),
    .D(\usb2uart.u_usb_cdc.u_sie.pid_q[0] ),
    .X(_2019_));
 sky130_fd_sc_hd__nor2_2 _2108_ (.A(\usb2uart.u_usb_cdc.out_err ),
    .B(_2019_),
    .Y(_2020_));
 sky130_fd_sc_hd__and3_1 _2109_ (.A(\usb2uart.u_usb_cdc.u_ctrl_endp.in_req_q ),
    .B(_2009_),
    .C(_2020_),
    .X(_2021_));
 sky130_fd_sc_hd__a21bo_1 _2110_ (.A1(_2011_),
    .A2(_2018_),
    .B1_N(_2021_),
    .X(_2022_));
 sky130_fd_sc_hd__buf_2 _2111_ (.A(\usb2uart.u_usb_cdc.u_ctrl_endp.byte_cnt_q[4] ),
    .X(_2023_));
 sky130_fd_sc_hd__clkinv_2 _2112_ (.A(\usb2uart.u_usb_cdc.u_ctrl_endp.byte_cnt_q[5] ),
    .Y(_2024_));
 sky130_fd_sc_hd__nand4b_2 _2113_ (.A_N(\usb2uart.u_usb_cdc.u_ctrl_endp.byte_cnt_q[2] ),
    .B(\usb2uart.u_usb_cdc.u_ctrl_endp.req_q[8] ),
    .C(\usb2uart.u_usb_cdc.u_ctrl_endp.byte_cnt_q[0] ),
    .D(\usb2uart.u_usb_cdc.u_ctrl_endp.byte_cnt_q[1] ),
    .Y(_2025_));
 sky130_fd_sc_hd__nor2_1 _2114_ (.A(\usb2uart.u_usb_cdc.u_ctrl_endp.byte_cnt_q[3] ),
    .B(_2025_),
    .Y(_2026_));
 sky130_fd_sc_hd__and4b_1 _2115_ (.A_N(_2023_),
    .B(_2024_),
    .C(\usb2uart.u_usb_cdc.u_ctrl_endp.byte_cnt_q[6] ),
    .D(_2026_),
    .X(_2027_));
 sky130_fd_sc_hd__xor2_1 _2116_ (.A(\usb2uart.u_usb_cdc.u_ctrl_endp.max_length_q[2] ),
    .B(\usb2uart.u_usb_cdc.u_ctrl_endp.byte_cnt_q[2] ),
    .X(_2028_));
 sky130_fd_sc_hd__xor2_1 _2117_ (.A(\usb2uart.u_usb_cdc.u_ctrl_endp.max_length_q[5] ),
    .B(\usb2uart.u_usb_cdc.u_ctrl_endp.byte_cnt_q[5] ),
    .X(_2029_));
 sky130_fd_sc_hd__xor2_1 _2118_ (.A(\usb2uart.u_usb_cdc.u_ctrl_endp.max_length_q[0] ),
    .B(\usb2uart.u_usb_cdc.u_ctrl_endp.byte_cnt_q[0] ),
    .X(_2030_));
 sky130_fd_sc_hd__xor2_1 _2119_ (.A(\usb2uart.u_usb_cdc.u_ctrl_endp.max_length_q[3] ),
    .B(\usb2uart.u_usb_cdc.u_ctrl_endp.byte_cnt_q[3] ),
    .X(_2031_));
 sky130_fd_sc_hd__or4_1 _2120_ (.A(_2028_),
    .B(_2029_),
    .C(_2030_),
    .D(_2031_),
    .X(_2032_));
 sky130_fd_sc_hd__or2_1 _2121_ (.A(\usb2uart.u_usb_cdc.u_ctrl_endp.max_length_q[4] ),
    .B(_2023_),
    .X(_2033_));
 sky130_fd_sc_hd__nand2_1 _2122_ (.A(\usb2uart.u_usb_cdc.u_ctrl_endp.max_length_q[4] ),
    .B(_2023_),
    .Y(_2034_));
 sky130_fd_sc_hd__or2_1 _2123_ (.A(\usb2uart.u_usb_cdc.u_ctrl_endp.max_length_q[1] ),
    .B(\usb2uart.u_usb_cdc.u_ctrl_endp.byte_cnt_q[1] ),
    .X(_2035_));
 sky130_fd_sc_hd__nand2_1 _2124_ (.A(\usb2uart.u_usb_cdc.u_ctrl_endp.max_length_q[1] ),
    .B(\usb2uart.u_usb_cdc.u_ctrl_endp.byte_cnt_q[1] ),
    .Y(_2036_));
 sky130_fd_sc_hd__xor2_1 _2125_ (.A(\usb2uart.u_usb_cdc.u_ctrl_endp.max_length_q[6] ),
    .B(\usb2uart.u_usb_cdc.u_ctrl_endp.byte_cnt_q[6] ),
    .X(_2037_));
 sky130_fd_sc_hd__a221o_1 _2126_ (.A1(_2033_),
    .A2(_2034_),
    .B1(_2035_),
    .B2(_2036_),
    .C1(_2037_),
    .X(_2038_));
 sky130_fd_sc_hd__and2b_1 _2127_ (.A_N(\usb2uart.u_usb_cdc.u_ctrl_endp.byte_cnt_q[0] ),
    .B(\usb2uart.u_usb_cdc.u_ctrl_endp.byte_cnt_q[1] ),
    .X(_2039_));
 sky130_fd_sc_hd__nor2_1 _2128_ (.A(\usb2uart.u_usb_cdc.u_ctrl_endp.byte_cnt_q[2] ),
    .B(\usb2uart.u_usb_cdc.u_ctrl_endp.byte_cnt_q[3] ),
    .Y(_2040_));
 sky130_fd_sc_hd__and4bb_1 _2129_ (.A_N(\usb2uart.u_usb_cdc.u_ctrl_endp.byte_cnt_q[5] ),
    .B_N(\usb2uart.u_usb_cdc.u_ctrl_endp.byte_cnt_q[6] ),
    .C(\usb2uart.u_usb_cdc.u_ctrl_endp.req_q[2] ),
    .D(_2023_),
    .X(_2041_));
 sky130_fd_sc_hd__and3_1 _2130_ (.A(_2039_),
    .B(_2040_),
    .C(_2041_),
    .X(_2042_));
 sky130_fd_sc_hd__o21ba_1 _2131_ (.A1(_2032_),
    .A2(_2038_),
    .B1_N(_2042_),
    .X(_2043_));
 sky130_fd_sc_hd__inv_2 _2132_ (.A(\usb2uart.u_usb_cdc.u_ctrl_endp.req_q[3] ),
    .Y(_2044_));
 sky130_fd_sc_hd__xnor2_2 _2133_ (.A(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.rx_valid_fq ),
    .B(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.rx_valid_fd ),
    .Y(_2045_));
 sky130_fd_sc_hd__or3b_1 _2134_ (.A(_2045_),
    .B(\usb2uart.u_usb_cdc.u_sie.rx_err ),
    .C_N(\usb2uart.u_usb_cdc.u_sie.phy_state_q[8] ),
    .X(_2046_));
 sky130_fd_sc_hd__o211a_1 _2135_ (.A1(_2044_),
    .A2(\usb2uart.u_usb_cdc.u_ctrl_endp.dev_state_qq[1] ),
    .B1(\usb2uart.u_usb_cdc.u_ctrl_endp.state_q[3] ),
    .C1(_2046_),
    .X(_2047_));
 sky130_fd_sc_hd__nand4b_2 _2136_ (.A_N(_2027_),
    .B(_2043_),
    .C(_2047_),
    .D(_2021_),
    .Y(_2048_));
 sky130_fd_sc_hd__and2_1 _2137_ (.A(\usb2uart.u_usb_cdc.endp[0] ),
    .B(_2007_),
    .X(_2049_));
 sky130_fd_sc_hd__nand2_1 _2138_ (.A(\usb2uart.u_usb_cdc.bulk_in_valid ),
    .B(_2049_),
    .Y(_2050_));
 sky130_fd_sc_hd__nand3_2 _2139_ (.A(_2022_),
    .B(_2048_),
    .C(_2050_),
    .Y(_2051_));
 sky130_fd_sc_hd__inv_2 _2140_ (.A(\usb2uart.u_usb_cdc.u_sie.in_byte_q[2] ),
    .Y(_2052_));
 sky130_fd_sc_hd__nand2_1 _2141_ (.A(\usb2uart.u_usb_cdc.u_sie.in_byte_q[1] ),
    .B(\usb2uart.u_usb_cdc.u_sie.in_byte_q[0] ),
    .Y(_2053_));
 sky130_fd_sc_hd__or3_2 _2142_ (.A(_2052_),
    .B(\usb2uart.u_usb_cdc.u_sie.in_byte_q[3] ),
    .C(_2053_),
    .X(_2054_));
 sky130_fd_sc_hd__nand2_2 _2143_ (.A(\usb2uart.u_usb_cdc.ctrl_stall ),
    .B(_2009_),
    .Y(_2055_));
 sky130_fd_sc_hd__and2_2 _2144_ (.A(\usb2uart.u_usb_cdc.u_sie.phy_state_q[1] ),
    .B(_2055_),
    .X(_2056_));
 sky130_fd_sc_hd__a21boi_2 _2145_ (.A1(_2048_),
    .A2(_2050_),
    .B1_N(_2022_),
    .Y(_2057_));
 sky130_fd_sc_hd__a32oi_4 _2146_ (.A1(\usb2uart.u_usb_cdc.u_sie.phy_state_q[7] ),
    .A2(_2051_),
    .A3(_2054_),
    .B1(_2056_),
    .B2(_2057_),
    .Y(_2058_));
 sky130_fd_sc_hd__nand2_1 _2147_ (.A(\usb2uart.u_usb_cdc.u_sie.u_phy_tx.stuffing_cnt_q[1] ),
    .B(\usb2uart.u_usb_cdc.u_sie.u_phy_tx.stuffing_cnt_q[2] ),
    .Y(_2059_));
 sky130_fd_sc_hd__or2_1 _2148_ (.A(\usb2uart.u_usb_cdc.u_sie.u_phy_tx.stuffing_cnt_q[0] ),
    .B(_2059_),
    .X(_2060_));
 sky130_fd_sc_hd__and3_1 _2149_ (.A(\usb2uart.u_usb_cdc.u_sie.u_phy_tx.clk_cnt_q[1] ),
    .B(\usb2uart.u_usb_cdc.u_sie.u_phy_tx.clk_cnt_q[0] ),
    .C(_2060_),
    .X(_2061_));
 sky130_fd_sc_hd__nand2_1 _2150_ (.A(\usb2uart.u_usb_cdc.u_sie.u_phy_tx.tx_valid_q ),
    .B(_2061_),
    .Y(_2062_));
 sky130_fd_sc_hd__or3_2 _2151_ (.A(\usb2uart.u_usb_cdc.u_sie.u_phy_tx.bit_cnt_q[2] ),
    .B(\usb2uart.u_usb_cdc.u_sie.u_phy_tx.bit_cnt_q[0] ),
    .C(\usb2uart.u_usb_cdc.u_sie.u_phy_tx.bit_cnt_q[1] ),
    .X(_2063_));
 sky130_fd_sc_hd__or4_4 _2152_ (.A(net6),
    .B(\usb2uart.u_usb_cdc.u_sie.u_phy_tx.tx_state_q[3] ),
    .C(_2062_),
    .D(_2063_),
    .X(_2064_));
 sky130_fd_sc_hd__and3b_1 _2153_ (.A_N(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.stuffing_cnt_q[0] ),
    .B(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.stuffing_cnt_q[1] ),
    .C(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.stuffing_cnt_q[2] ),
    .X(_2065_));
 sky130_fd_sc_hd__or2b_1 _2154_ (.A(_2065_),
    .B_N(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.data_q[0] ),
    .X(_2066_));
 sky130_fd_sc_hd__inv_2 _2155_ (.A(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.nrzi_q[3] ),
    .Y(_2067_));
 sky130_fd_sc_hd__a31o_1 _2156_ (.A1(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.nrzi_q[2] ),
    .A2(_2067_),
    .A3(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.rx_state_q[4] ),
    .B1(\usb2uart.u_usb_cdc.u_sie.rx_err ),
    .X(_2068_));
 sky130_fd_sc_hd__inv_2 _2157_ (.A(_2068_),
    .Y(_2069_));
 sky130_fd_sc_hd__nand2b_2 _2158_ (.A_N(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.clk_cnt_q[1] ),
    .B(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.clk_cnt_q[0] ),
    .Y(_2070_));
 sky130_fd_sc_hd__a21o_1 _2159_ (.A1(_2066_),
    .A2(_2069_),
    .B1(_2070_),
    .X(_2071_));
 sky130_fd_sc_hd__and3_1 _2160_ (.A(\usb2uart.u_usb_cdc.u_sie.delay_cnt_q[1] ),
    .B(\usb2uart.u_usb_cdc.u_sie.delay_cnt_q[0] ),
    .C(\usb2uart.u_usb_cdc.u_sie.delay_cnt_q[2] ),
    .X(_2072_));
 sky130_fd_sc_hd__and2_1 _2161_ (.A(\usb2uart.u_usb_cdc.u_sie.delay_cnt_q[3] ),
    .B(_2072_),
    .X(_2073_));
 sky130_fd_sc_hd__nand2_1 _2162_ (.A(\usb2uart.u_usb_cdc.u_sie.delay_cnt_q[4] ),
    .B(_2073_),
    .Y(_2074_));
 sky130_fd_sc_hd__clkbuf_2 _2163_ (.A(\usb2uart.u_usb_cdc.out_err ),
    .X(_2075_));
 sky130_fd_sc_hd__nor2_1 _2164_ (.A(_2075_),
    .B(\usb2uart.u_usb_cdc.u_sie.out_eop_q ),
    .Y(_2076_));
 sky130_fd_sc_hd__o22a_1 _2165_ (.A1(_2046_),
    .A2(_2071_),
    .B1(_2074_),
    .B2(_2076_),
    .X(_2077_));
 sky130_fd_sc_hd__o31ai_4 _2166_ (.A1(\usb2uart.u_usb_cdc.u_sie.rx_err ),
    .A2(_2058_),
    .A3(_2064_),
    .B1(_2077_),
    .Y(_2078_));
 sky130_fd_sc_hd__and3_1 _2167_ (.A(_2006_),
    .B(_2009_),
    .C(_2078_),
    .X(_2079_));
 sky130_fd_sc_hd__buf_2 _2168_ (.A(_2079_),
    .X(_2080_));
 sky130_fd_sc_hd__or2_2 _2169_ (.A(_2075_),
    .B(_2019_),
    .X(_2081_));
 sky130_fd_sc_hd__nor2_2 _2170_ (.A(_2012_),
    .B(_2081_),
    .Y(_2082_));
 sky130_fd_sc_hd__clkbuf_4 _2171_ (.A(\usb2uart.u_usb_cdc.u_ctrl_endp.byte_cnt_q[0] ),
    .X(_2083_));
 sky130_fd_sc_hd__clkinv_2 _2172_ (.A(_2083_),
    .Y(_2084_));
 sky130_fd_sc_hd__buf_2 _2173_ (.A(\usb2uart.u_usb_cdc.u_ctrl_endp.byte_cnt_q[1] ),
    .X(_0450_));
 sky130_fd_sc_hd__nor2_1 _2174_ (.A(_2084_),
    .B(_0450_),
    .Y(_0451_));
 sky130_fd_sc_hd__buf_2 _2175_ (.A(\usb2uart.u_usb_cdc.u_ctrl_endp.byte_cnt_q[2] ),
    .X(_0452_));
 sky130_fd_sc_hd__clkbuf_4 _2176_ (.A(\usb2uart.u_usb_cdc.u_ctrl_endp.byte_cnt_q[3] ),
    .X(_0453_));
 sky130_fd_sc_hd__buf_2 _2177_ (.A(\usb2uart.u_usb_cdc.u_ctrl_endp.byte_cnt_q[5] ),
    .X(_0454_));
 sky130_fd_sc_hd__or3_1 _2178_ (.A(_2023_),
    .B(_0454_),
    .C(\usb2uart.u_usb_cdc.u_ctrl_endp.byte_cnt_q[6] ),
    .X(_0455_));
 sky130_fd_sc_hd__or2_1 _2179_ (.A(_0453_),
    .B(_0455_),
    .X(_0456_));
 sky130_fd_sc_hd__nor2_1 _2180_ (.A(_0452_),
    .B(_0456_),
    .Y(_0457_));
 sky130_fd_sc_hd__and2_1 _2181_ (.A(_0451_),
    .B(_0457_),
    .X(_0458_));
 sky130_fd_sc_hd__and3_1 _2182_ (.A(\usb2uart.u_usb_cdc.u_ctrl_endp.req_q[0] ),
    .B(_2082_),
    .C(_0458_),
    .X(_0459_));
 sky130_fd_sc_hd__and3_1 _2183_ (.A(_2002_),
    .B(_2080_),
    .C(_0459_),
    .X(_0460_));
 sky130_fd_sc_hd__clkbuf_4 _2184_ (.A(\usb2uart.u_usb_cdc.u_ctrl_endp.in_dir_q ),
    .X(_0461_));
 sky130_fd_sc_hd__or2_1 _2185_ (.A(\usb2uart.u_usb_cdc.u_ctrl_endp.rec_q[0] ),
    .B(\usb2uart.u_usb_cdc.u_ctrl_endp.rec_q[1] ),
    .X(_0462_));
 sky130_fd_sc_hd__nor2_1 _2186_ (.A(_0461_),
    .B(_0462_),
    .Y(_0463_));
 sky130_fd_sc_hd__inv_2 _2187_ (.A(\usb2uart.u_usb_cdc.out_data[0] ),
    .Y(_0464_));
 sky130_fd_sc_hd__clkbuf_4 _2188_ (.A(\usb2uart.u_usb_cdc.out_data[1] ),
    .X(_0465_));
 sky130_fd_sc_hd__clkbuf_4 _2189_ (.A(\usb2uart.u_usb_cdc.out_data[6] ),
    .X(_0466_));
 sky130_fd_sc_hd__or3_1 _2190_ (.A(\usb2uart.u_usb_cdc.out_data[4] ),
    .B(\usb2uart.u_usb_cdc.out_data[5] ),
    .C(_0466_),
    .X(_0467_));
 sky130_fd_sc_hd__or2_2 _2191_ (.A(\usb2uart.u_usb_cdc.out_data[7] ),
    .B(_0467_),
    .X(_0468_));
 sky130_fd_sc_hd__inv_2 _2192_ (.A(\usb2uart.u_usb_cdc.out_data[3] ),
    .Y(_0469_));
 sky130_fd_sc_hd__nand2_1 _2193_ (.A(\usb2uart.u_usb_cdc.out_data[2] ),
    .B(_0469_),
    .Y(_0470_));
 sky130_fd_sc_hd__or4_1 _2194_ (.A(_0464_),
    .B(_0465_),
    .C(_0468_),
    .D(_0470_),
    .X(_0471_));
 sky130_fd_sc_hd__inv_2 _2195_ (.A(_0471_),
    .Y(_0472_));
 sky130_fd_sc_hd__buf_2 _2196_ (.A(\usb2uart.u_usb_cdc.u_ctrl_endp.state_q[1] ),
    .X(_0473_));
 sky130_fd_sc_hd__nand2_2 _2197_ (.A(_0473_),
    .B(_2020_),
    .Y(_0474_));
 sky130_fd_sc_hd__nor2_1 _2198_ (.A(_0453_),
    .B(_0455_),
    .Y(_0475_));
 sky130_fd_sc_hd__nand2_1 _2199_ (.A(\usb2uart.u_usb_cdc.u_ctrl_endp.byte_cnt_q[2] ),
    .B(_0475_),
    .Y(_0476_));
 sky130_fd_sc_hd__clkinv_2 _2200_ (.A(_0450_),
    .Y(_0477_));
 sky130_fd_sc_hd__nand2_2 _2201_ (.A(_2083_),
    .B(_0477_),
    .Y(_0478_));
 sky130_fd_sc_hd__nor3_2 _2202_ (.A(_0474_),
    .B(_0476_),
    .C(_0478_),
    .Y(_0479_));
 sky130_fd_sc_hd__nor2_1 _2203_ (.A(_2084_),
    .B(_0477_),
    .Y(_0480_));
 sky130_fd_sc_hd__and3_1 _2204_ (.A(_0480_),
    .B(_2082_),
    .C(_0457_),
    .X(_0481_));
 sky130_fd_sc_hd__clkbuf_4 _2205_ (.A(\usb2uart.u_usb_cdc.out_data[0] ),
    .X(_0482_));
 sky130_fd_sc_hd__or2_2 _2206_ (.A(\usb2uart.u_usb_cdc.out_data[2] ),
    .B(\usb2uart.u_usb_cdc.out_data[3] ),
    .X(_0483_));
 sky130_fd_sc_hd__or3_4 _2207_ (.A(\usb2uart.u_usb_cdc.out_data[1] ),
    .B(_0483_),
    .C(_0468_),
    .X(_0484_));
 sky130_fd_sc_hd__nor2_4 _2208_ (.A(_0482_),
    .B(_0484_),
    .Y(_0485_));
 sky130_fd_sc_hd__o211a_1 _2209_ (.A1(_0479_),
    .A2(_0481_),
    .B1(_2080_),
    .C1(_0485_),
    .X(_0486_));
 sky130_fd_sc_hd__clkbuf_4 _2210_ (.A(_2046_),
    .X(_0487_));
 sky130_fd_sc_hd__nand2_1 _2211_ (.A(_2009_),
    .B(_2078_),
    .Y(_0488_));
 sky130_fd_sc_hd__nand2_1 _2212_ (.A(_2039_),
    .B(_0457_),
    .Y(_0489_));
 sky130_fd_sc_hd__or4_2 _2213_ (.A(_0487_),
    .B(_0488_),
    .C(_0474_),
    .D(_0489_),
    .X(_0490_));
 sky130_fd_sc_hd__nor2_1 _2214_ (.A(\usb2uart.u_usb_cdc.out_data[7] ),
    .B(_0490_),
    .Y(_0491_));
 sky130_fd_sc_hd__nor2_2 _2215_ (.A(_2083_),
    .B(\usb2uart.u_usb_cdc.u_ctrl_endp.byte_cnt_q[1] ),
    .Y(_0492_));
 sky130_fd_sc_hd__and2_1 _2216_ (.A(_0452_),
    .B(_0492_),
    .X(_0493_));
 sky130_fd_sc_hd__inv_2 _2217_ (.A(_0493_),
    .Y(_0494_));
 sky130_fd_sc_hd__nor2_2 _2218_ (.A(_0456_),
    .B(_0494_),
    .Y(_0495_));
 sky130_fd_sc_hd__and4_1 _2219_ (.A(_2006_),
    .B(_0485_),
    .C(_2082_),
    .D(_0495_),
    .X(_0496_));
 sky130_fd_sc_hd__nor2_1 _2220_ (.A(_2012_),
    .B(_2006_),
    .Y(_0497_));
 sky130_fd_sc_hd__or3_2 _2221_ (.A(\usb2uart.u_usb_cdc.u_ctrl_endp.state_q[3] ),
    .B(\usb2uart.u_usb_cdc.ctrl_stall ),
    .C(\usb2uart.u_usb_cdc.u_ctrl_endp.state_q[0] ),
    .X(_0498_));
 sky130_fd_sc_hd__or2_1 _2222_ (.A(_0497_),
    .B(_0498_),
    .X(_0499_));
 sky130_fd_sc_hd__or4_1 _2223_ (.A(_2075_),
    .B(_2019_),
    .C(_0488_),
    .D(_0499_),
    .X(_0500_));
 sky130_fd_sc_hd__and3_1 _2224_ (.A(_2083_),
    .B(\usb2uart.u_usb_cdc.u_ctrl_endp.byte_cnt_q[1] ),
    .C(\usb2uart.u_usb_cdc.u_ctrl_endp.byte_cnt_q[2] ),
    .X(_0501_));
 sky130_fd_sc_hd__buf_2 _2225_ (.A(_0501_),
    .X(_0502_));
 sky130_fd_sc_hd__nand2_1 _2226_ (.A(_0475_),
    .B(_0502_),
    .Y(_0503_));
 sky130_fd_sc_hd__nor2_1 _2227_ (.A(_0474_),
    .B(_0503_),
    .Y(_0504_));
 sky130_fd_sc_hd__or2_1 _2228_ (.A(\usb2uart.u_usb_cdc.u_ctrl_endp.req_q[3] ),
    .B(\usb2uart.u_usb_cdc.u_ctrl_endp.req_q[5] ),
    .X(_0505_));
 sky130_fd_sc_hd__nand2_1 _2229_ (.A(_2084_),
    .B(_0450_),
    .Y(_0506_));
 sky130_fd_sc_hd__or3_1 _2230_ (.A(_0506_),
    .B(_0474_),
    .C(_0476_),
    .X(_0507_));
 sky130_fd_sc_hd__nor2_1 _2231_ (.A(_0505_),
    .B(_0507_),
    .Y(_0508_));
 sky130_fd_sc_hd__o211a_1 _2232_ (.A1(_0504_),
    .A2(_0508_),
    .B1(_2079_),
    .C1(_0485_),
    .X(_0509_));
 sky130_fd_sc_hd__or3_1 _2233_ (.A(_0496_),
    .B(_0500_),
    .C(_0509_),
    .X(_0510_));
 sky130_fd_sc_hd__and3_1 _2234_ (.A(_2079_),
    .B(_2082_),
    .C(_0456_),
    .X(_0511_));
 sky130_fd_sc_hd__o41a_1 _2235_ (.A1(_0486_),
    .A2(_0491_),
    .A3(_0510_),
    .A4(_0511_),
    .B1(\usb2uart.u_usb_cdc.u_ctrl_endp.req_q[1] ),
    .X(_0512_));
 sky130_fd_sc_hd__a31o_1 _2236_ (.A1(_0460_),
    .A2(_0463_),
    .A3(_0472_),
    .B1(_0512_),
    .X(_0004_));
 sky130_fd_sc_hd__and2_1 _2237_ (.A(_2071_),
    .B(_2064_),
    .X(_0513_));
 sky130_fd_sc_hd__clkbuf_4 _2238_ (.A(_0513_),
    .X(_0514_));
 sky130_fd_sc_hd__clkbuf_4 _2239_ (.A(_0514_),
    .X(_0515_));
 sky130_fd_sc_hd__nand2_4 _2240_ (.A(_2071_),
    .B(_2064_),
    .Y(_0516_));
 sky130_fd_sc_hd__clkbuf_4 _2241_ (.A(\usb2uart.u_usb_cdc.u_sie.data_q[0] ),
    .X(_0517_));
 sky130_fd_sc_hd__clkbuf_4 _2242_ (.A(\usb2uart.u_usb_cdc.u_sie.phy_state_q[6] ),
    .X(_0518_));
 sky130_fd_sc_hd__buf_4 _2243_ (.A(\usb2uart.u_usb_cdc.u_sie.data_q[3] ),
    .X(_0519_));
 sky130_fd_sc_hd__xnor2_1 _2244_ (.A(\usb2uart.u_usb_cdc.u_sie.data_q[7] ),
    .B(_0519_),
    .Y(_0520_));
 sky130_fd_sc_hd__clkbuf_4 _2245_ (.A(\usb2uart.u_usb_cdc.u_sie.data_q[1] ),
    .X(_0521_));
 sky130_fd_sc_hd__a2bb2o_1 _2246_ (.A1_N(_0521_),
    .A2_N(\usb2uart.u_usb_cdc.u_sie.data_q[5] ),
    .B1(\usb2uart.u_usb_cdc.u_sie.data_q[4] ),
    .B2(\usb2uart.u_usb_cdc.u_sie.data_q[0] ),
    .X(_0522_));
 sky130_fd_sc_hd__a2bb2o_1 _2247_ (.A1_N(\usb2uart.u_usb_cdc.u_sie.data_q[0] ),
    .A2_N(\usb2uart.u_usb_cdc.u_sie.data_q[4] ),
    .B1(\usb2uart.u_usb_cdc.u_sie.data_q[5] ),
    .B2(_0521_),
    .X(_0523_));
 sky130_fd_sc_hd__or3_1 _2248_ (.A(_0520_),
    .B(_0522_),
    .C(_0523_),
    .X(_0524_));
 sky130_fd_sc_hd__or3b_1 _2249_ (.A(_0524_),
    .B(\usb2uart.u_usb_cdc.u_sie.data_q[6] ),
    .C_N(\usb2uart.u_usb_cdc.u_sie.data_q[2] ),
    .X(_0525_));
 sky130_fd_sc_hd__or3b_1 _2250_ (.A(\usb2uart.u_usb_cdc.u_sie.data_q[2] ),
    .B(_0524_),
    .C_N(\usb2uart.u_usb_cdc.u_sie.data_q[6] ),
    .X(_0526_));
 sky130_fd_sc_hd__nand2_2 _2251_ (.A(_0525_),
    .B(_0526_),
    .Y(_0527_));
 sky130_fd_sc_hd__and4_1 _2252_ (.A(_2003_),
    .B(_0517_),
    .C(_0518_),
    .D(_0527_),
    .X(_0528_));
 sky130_fd_sc_hd__and3_1 _2253_ (.A(_2004_),
    .B(_0516_),
    .C(_0528_),
    .X(_0529_));
 sky130_fd_sc_hd__clkinv_2 _2254_ (.A(\usb2uart.u_usb_cdc.u_sie.data_q[1] ),
    .Y(_0530_));
 sky130_fd_sc_hd__a22o_1 _2255_ (.A1(\usb2uart.u_usb_cdc.u_sie.phy_state_q[3] ),
    .A2(_0515_),
    .B1(_0529_),
    .B2(_0530_),
    .X(_0022_));
 sky130_fd_sc_hd__inv_2 _2256_ (.A(\usb2uart.u_usb_cdc.u_sie.pid_q[3] ),
    .Y(_0531_));
 sky130_fd_sc_hd__inv_2 _2257_ (.A(\usb2uart.u_usb_cdc.u_sie.pid_q[2] ),
    .Y(_0532_));
 sky130_fd_sc_hd__or2b_1 _2258_ (.A(\usb2uart.u_usb_cdc.u_sie.pid_q[1] ),
    .B_N(\usb2uart.u_usb_cdc.u_sie.pid_q[0] ),
    .X(_0533_));
 sky130_fd_sc_hd__or3_2 _2259_ (.A(_0531_),
    .B(_0532_),
    .C(_0533_),
    .X(_0534_));
 sky130_fd_sc_hd__or3_1 _2260_ (.A(\usb2uart.u_usb_cdc.u_sie.pid_q[3] ),
    .B(\usb2uart.u_usb_cdc.u_sie.pid_q[2] ),
    .C(_0533_),
    .X(_0535_));
 sky130_fd_sc_hd__inv_2 _2261_ (.A(\usb2uart.u_usb_cdc.addr[4] ),
    .Y(_0536_));
 sky130_fd_sc_hd__inv_2 _2262_ (.A(\usb2uart.u_usb_cdc.u_sie.addr_q[5] ),
    .Y(_0537_));
 sky130_fd_sc_hd__xor2_1 _2263_ (.A(\usb2uart.u_usb_cdc.u_sie.addr_q[1] ),
    .B(\usb2uart.u_usb_cdc.addr[1] ),
    .X(_0538_));
 sky130_fd_sc_hd__a221o_1 _2264_ (.A1(\usb2uart.u_usb_cdc.u_sie.addr_q[4] ),
    .A2(_0536_),
    .B1(_0537_),
    .B2(\usb2uart.u_usb_cdc.addr[5] ),
    .C1(_0538_),
    .X(_0539_));
 sky130_fd_sc_hd__inv_2 _2265_ (.A(\usb2uart.u_usb_cdc.u_sie.addr_q[0] ),
    .Y(_0540_));
 sky130_fd_sc_hd__nand2_1 _2266_ (.A(\usb2uart.u_usb_cdc.u_sie.addr_q[6] ),
    .B(\usb2uart.u_usb_cdc.addr[6] ),
    .Y(_0541_));
 sky130_fd_sc_hd__or2_1 _2267_ (.A(\usb2uart.u_usb_cdc.u_sie.addr_q[6] ),
    .B(\usb2uart.u_usb_cdc.addr[6] ),
    .X(_0542_));
 sky130_fd_sc_hd__a221o_1 _2268_ (.A1(_0540_),
    .A2(\usb2uart.u_usb_cdc.addr[0] ),
    .B1(_0541_),
    .B2(_0542_),
    .C1(\usb2uart.u_usb_cdc.u_sie.data_q[2] ),
    .X(_0543_));
 sky130_fd_sc_hd__inv_2 _2269_ (.A(\usb2uart.u_usb_cdc.addr[2] ),
    .Y(_0544_));
 sky130_fd_sc_hd__o2bb2a_1 _2270_ (.A1_N(\usb2uart.u_usb_cdc.u_sie.addr_q[2] ),
    .A2_N(_0544_),
    .B1(_0537_),
    .B2(\usb2uart.u_usb_cdc.addr[5] ),
    .X(_0545_));
 sky130_fd_sc_hd__inv_2 _2271_ (.A(\usb2uart.u_usb_cdc.u_sie.addr_q[3] ),
    .Y(_0546_));
 sky130_fd_sc_hd__inv_2 _2272_ (.A(\usb2uart.u_usb_cdc.addr[3] ),
    .Y(_0547_));
 sky130_fd_sc_hd__o22a_1 _2273_ (.A1(\usb2uart.u_usb_cdc.u_sie.addr_q[3] ),
    .A2(_0547_),
    .B1(\usb2uart.u_usb_cdc.u_sie.addr_q[4] ),
    .B2(_0536_),
    .X(_0548_));
 sky130_fd_sc_hd__o221a_1 _2274_ (.A1(_0540_),
    .A2(\usb2uart.u_usb_cdc.addr[0] ),
    .B1(_0546_),
    .B2(\usb2uart.u_usb_cdc.addr[3] ),
    .C1(_0548_),
    .X(_0549_));
 sky130_fd_sc_hd__o211a_1 _2275_ (.A1(\usb2uart.u_usb_cdc.u_sie.addr_q[2] ),
    .A2(_0544_),
    .B1(_0545_),
    .C1(_0549_),
    .X(_0550_));
 sky130_fd_sc_hd__or3b_2 _2276_ (.A(_0539_),
    .B(_0543_),
    .C_N(_0550_),
    .X(_0551_));
 sky130_fd_sc_hd__a21oi_1 _2277_ (.A1(_0534_),
    .A2(_0535_),
    .B1(_0551_),
    .Y(_0552_));
 sky130_fd_sc_hd__a32o_1 _2278_ (.A1(_0521_),
    .A2(_0529_),
    .A3(_0552_),
    .B1(\usb2uart.u_usb_cdc.u_sie.phy_state_q[2] ),
    .B2(_0514_),
    .X(_0021_));
 sky130_fd_sc_hd__clkbuf_4 _2279_ (.A(\usb2uart.u_usb_cdc.u_sie.phy_state_q[1] ),
    .X(_0553_));
 sky130_fd_sc_hd__inv_2 _2280_ (.A(\usb2uart.u_usb_cdc.u_sie.data_q[7] ),
    .Y(_0554_));
 sky130_fd_sc_hd__xor2_1 _2281_ (.A(\usb2uart.u_usb_cdc.out_data[1] ),
    .B(\usb2uart.u_usb_cdc.out_data[4] ),
    .X(_0555_));
 sky130_fd_sc_hd__xnor2_1 _2282_ (.A(\usb2uart.u_usb_cdc.out_data[2] ),
    .B(\usb2uart.u_usb_cdc.out_data[7] ),
    .Y(_0556_));
 sky130_fd_sc_hd__xnor2_1 _2283_ (.A(_0555_),
    .B(_0556_),
    .Y(_0557_));
 sky130_fd_sc_hd__xnor2_1 _2284_ (.A(\usb2uart.u_usb_cdc.out_data[2] ),
    .B(\usb2uart.u_usb_cdc.out_data[5] ),
    .Y(_0558_));
 sky130_fd_sc_hd__xnor2_1 _2285_ (.A(\usb2uart.u_usb_cdc.out_data[0] ),
    .B(_0558_),
    .Y(_0559_));
 sky130_fd_sc_hd__xnor2_1 _2286_ (.A(\usb2uart.u_usb_cdc.u_sie.data_q[2] ),
    .B(_0559_),
    .Y(_0560_));
 sky130_fd_sc_hd__xnor2_1 _2287_ (.A(_0557_),
    .B(_0560_),
    .Y(_0561_));
 sky130_fd_sc_hd__xor2_1 _2288_ (.A(\usb2uart.u_usb_cdc.out_data[0] ),
    .B(\usb2uart.u_usb_cdc.out_data[3] ),
    .X(_0562_));
 sky130_fd_sc_hd__xnor2_1 _2289_ (.A(_0530_),
    .B(_0562_),
    .Y(_0563_));
 sky130_fd_sc_hd__xor2_1 _2290_ (.A(\usb2uart.u_usb_cdc.out_data[4] ),
    .B(_0466_),
    .X(_0564_));
 sky130_fd_sc_hd__xnor2_1 _2291_ (.A(_0563_),
    .B(_0564_),
    .Y(_0565_));
 sky130_fd_sc_hd__xnor2_1 _2292_ (.A(\usb2uart.u_usb_cdc.u_sie.data_q[4] ),
    .B(_0557_),
    .Y(_0566_));
 sky130_fd_sc_hd__xor2_1 _2293_ (.A(\usb2uart.u_usb_cdc.out_data[1] ),
    .B(_0466_),
    .X(_0567_));
 sky130_fd_sc_hd__xnor2_1 _2294_ (.A(_0519_),
    .B(_0567_),
    .Y(_0568_));
 sky130_fd_sc_hd__xor2_1 _2295_ (.A(_0517_),
    .B(_0559_),
    .X(_0569_));
 sky130_fd_sc_hd__o2bb2a_1 _2296_ (.A1_N(_0565_),
    .A2_N(_0566_),
    .B1(_0568_),
    .B2(_0569_),
    .X(_0570_));
 sky130_fd_sc_hd__mux2_1 _2297_ (.A0(_0565_),
    .A1(_0566_),
    .S(\usb2uart.u_usb_cdc.u_sie.data_q[6] ),
    .X(_0571_));
 sky130_fd_sc_hd__o211ai_1 _2298_ (.A1(_0554_),
    .A2(_0561_),
    .B1(_0570_),
    .C1(_0571_),
    .Y(_0572_));
 sky130_fd_sc_hd__xnor2_1 _2299_ (.A(\usb2uart.u_usb_cdc.u_sie.data_q[5] ),
    .B(_0562_),
    .Y(_0573_));
 sky130_fd_sc_hd__xnor2_1 _2300_ (.A(_0561_),
    .B(_0573_),
    .Y(_0574_));
 sky130_fd_sc_hd__mux2_1 _2301_ (.A0(_0569_),
    .A1(_0568_),
    .S(_0574_),
    .X(_0575_));
 sky130_fd_sc_hd__a211o_1 _2302_ (.A1(_0554_),
    .A2(_0561_),
    .B1(_0572_),
    .C1(_0575_),
    .X(_0576_));
 sky130_fd_sc_hd__xor2_1 _2303_ (.A(_0466_),
    .B(\usb2uart.u_usb_cdc.addr[6] ),
    .X(_0577_));
 sky130_fd_sc_hd__xor2_1 _2304_ (.A(\usb2uart.u_usb_cdc.out_data[1] ),
    .B(\usb2uart.u_usb_cdc.addr[1] ),
    .X(_0578_));
 sky130_fd_sc_hd__a221o_1 _2305_ (.A1(\usb2uart.u_usb_cdc.out_data[2] ),
    .A2(_0544_),
    .B1(_0547_),
    .B2(\usb2uart.u_usb_cdc.out_data[3] ),
    .C1(_0578_),
    .X(_0579_));
 sky130_fd_sc_hd__inv_2 _2306_ (.A(\usb2uart.u_usb_cdc.addr[0] ),
    .Y(_0580_));
 sky130_fd_sc_hd__xor2_1 _2307_ (.A(\usb2uart.u_usb_cdc.out_data[4] ),
    .B(\usb2uart.u_usb_cdc.addr[4] ),
    .X(_0581_));
 sky130_fd_sc_hd__a221o_1 _2308_ (.A1(_0482_),
    .A2(_0580_),
    .B1(\usb2uart.u_usb_cdc.addr[3] ),
    .B2(_0469_),
    .C1(_0581_),
    .X(_0582_));
 sky130_fd_sc_hd__xnor2_1 _2309_ (.A(\usb2uart.u_usb_cdc.out_data[5] ),
    .B(\usb2uart.u_usb_cdc.addr[5] ),
    .Y(_0583_));
 sky130_fd_sc_hd__o221a_1 _2310_ (.A1(_0482_),
    .A2(_0580_),
    .B1(_0544_),
    .B2(\usb2uart.u_usb_cdc.out_data[2] ),
    .C1(_0583_),
    .X(_0584_));
 sky130_fd_sc_hd__or4b_2 _2311_ (.A(_0577_),
    .B(_0579_),
    .C(_0582_),
    .D_N(_0584_),
    .X(_0585_));
 sky130_fd_sc_hd__or4_1 _2312_ (.A(_0531_),
    .B(\usb2uart.u_usb_cdc.u_sie.pid_q[2] ),
    .C(_0533_),
    .D(_0585_),
    .X(_0586_));
 sky130_fd_sc_hd__nor2_1 _2313_ (.A(_0576_),
    .B(_0586_),
    .Y(_0587_));
 sky130_fd_sc_hd__buf_2 _2314_ (.A(_2045_),
    .X(_0588_));
 sky130_fd_sc_hd__clkbuf_4 _2315_ (.A(\usb2uart.u_usb_cdc.u_sie.rx_err ),
    .X(_0589_));
 sky130_fd_sc_hd__nor2_1 _2316_ (.A(_0589_),
    .B(_0514_),
    .Y(_0590_));
 sky130_fd_sc_hd__clkbuf_4 _2317_ (.A(_0590_),
    .X(_0591_));
 sky130_fd_sc_hd__and3_1 _2318_ (.A(\usb2uart.u_usb_cdc.u_sie.phy_state_q[9] ),
    .B(_0588_),
    .C(_0591_),
    .X(_0592_));
 sky130_fd_sc_hd__a22o_1 _2319_ (.A1(_0553_),
    .A2(_0515_),
    .B1(_0587_),
    .B2(_0592_),
    .X(_0020_));
 sky130_fd_sc_hd__inv_2 _2320_ (.A(\usb2uart.u_usb_cdc.u_sie.phy_state_q[9] ),
    .Y(_0593_));
 sky130_fd_sc_hd__nand2_1 _2321_ (.A(_0517_),
    .B(_0527_),
    .Y(_0594_));
 sky130_fd_sc_hd__nand2_1 _2322_ (.A(_0518_),
    .B(_0594_),
    .Y(_0595_));
 sky130_fd_sc_hd__o21ai_1 _2323_ (.A1(_0593_),
    .A2(_0587_),
    .B1(_0595_),
    .Y(_0596_));
 sky130_fd_sc_hd__clkbuf_4 _2324_ (.A(\usb2uart.u_usb_cdc.u_sie.phy_state_q[8] ),
    .X(_0597_));
 sky130_fd_sc_hd__xor2_1 _2325_ (.A(\usb2uart.u_usb_cdc.u_sie.data_q[7] ),
    .B(\usb2uart.u_usb_cdc.u_sie.crc16_q[8] ),
    .X(_0598_));
 sky130_fd_sc_hd__xnor2_2 _2326_ (.A(\usb2uart.u_usb_cdc.u_sie.data_q[2] ),
    .B(\usb2uart.u_usb_cdc.u_sie.crc16_q[13] ),
    .Y(_0599_));
 sky130_fd_sc_hd__xor2_2 _2327_ (.A(_0519_),
    .B(\usb2uart.u_usb_cdc.u_sie.crc16_q[12] ),
    .X(_0600_));
 sky130_fd_sc_hd__xnor2_2 _2328_ (.A(_0599_),
    .B(_0600_),
    .Y(_0601_));
 sky130_fd_sc_hd__xnor2_2 _2329_ (.A(\usb2uart.u_usb_cdc.u_sie.data_q[6] ),
    .B(\usb2uart.u_usb_cdc.u_sie.crc16_q[9] ),
    .Y(_0602_));
 sky130_fd_sc_hd__xnor2_1 _2330_ (.A(_0601_),
    .B(_0602_),
    .Y(_0603_));
 sky130_fd_sc_hd__xnor2_2 _2331_ (.A(\usb2uart.u_usb_cdc.u_sie.data_q[5] ),
    .B(\usb2uart.u_usb_cdc.u_sie.crc16_q[10] ),
    .Y(_0604_));
 sky130_fd_sc_hd__xor2_2 _2332_ (.A(\usb2uart.u_usb_cdc.u_sie.data_q[4] ),
    .B(\usb2uart.u_usb_cdc.u_sie.crc16_q[11] ),
    .X(_0605_));
 sky130_fd_sc_hd__xnor2_2 _2333_ (.A(_0604_),
    .B(_0605_),
    .Y(_0606_));
 sky130_fd_sc_hd__xor2_2 _2334_ (.A(\usb2uart.u_usb_cdc.u_sie.data_q[1] ),
    .B(\usb2uart.u_usb_cdc.u_sie.crc16_q[14] ),
    .X(_0607_));
 sky130_fd_sc_hd__xor2_2 _2335_ (.A(\usb2uart.u_usb_cdc.u_sie.data_q[0] ),
    .B(\usb2uart.u_usb_cdc.u_sie.crc16_q[15] ),
    .X(_0608_));
 sky130_fd_sc_hd__xor2_2 _2336_ (.A(_0607_),
    .B(_0608_),
    .X(_0609_));
 sky130_fd_sc_hd__xnor2_1 _2337_ (.A(_0606_),
    .B(_0609_),
    .Y(_0610_));
 sky130_fd_sc_hd__xnor2_1 _2338_ (.A(_0603_),
    .B(_0610_),
    .Y(_0611_));
 sky130_fd_sc_hd__inv_2 _2339_ (.A(_0611_),
    .Y(_0612_));
 sky130_fd_sc_hd__nand2_1 _2340_ (.A(_0598_),
    .B(_0612_),
    .Y(_0613_));
 sky130_fd_sc_hd__xor2_1 _2341_ (.A(\usb2uart.u_usb_cdc.u_sie.crc16_q[0] ),
    .B(_0609_),
    .X(_0614_));
 sky130_fd_sc_hd__xor2_1 _2342_ (.A(_0605_),
    .B(_0600_),
    .X(_0615_));
 sky130_fd_sc_hd__or3_1 _2343_ (.A(\usb2uart.u_usb_cdc.u_sie.crc16_q[5] ),
    .B(\usb2uart.u_usb_cdc.u_sie.crc16_q[4] ),
    .C(\usb2uart.u_usb_cdc.u_sie.crc16_q[6] ),
    .X(_0616_));
 sky130_fd_sc_hd__or3_1 _2344_ (.A(\usb2uart.u_usb_cdc.u_sie.crc16_q[3] ),
    .B(\usb2uart.u_usb_cdc.u_sie.crc16_q[2] ),
    .C(_0616_),
    .X(_0617_));
 sky130_fd_sc_hd__or3_1 _2345_ (.A(_0606_),
    .B(_0601_),
    .C(_0617_),
    .X(_0618_));
 sky130_fd_sc_hd__inv_2 _2346_ (.A(\usb2uart.u_usb_cdc.u_sie.crc16_q[1] ),
    .Y(_0619_));
 sky130_fd_sc_hd__xnor2_1 _2347_ (.A(_0619_),
    .B(_0608_),
    .Y(_0620_));
 sky130_fd_sc_hd__xnor2_1 _2348_ (.A(_0599_),
    .B(_0607_),
    .Y(_0621_));
 sky130_fd_sc_hd__xnor2_1 _2349_ (.A(_0598_),
    .B(_0602_),
    .Y(_0622_));
 sky130_fd_sc_hd__xor2_1 _2350_ (.A(_0604_),
    .B(_0602_),
    .X(_0623_));
 sky130_fd_sc_hd__or4bb_1 _2351_ (.A(_0620_),
    .B(_0621_),
    .C_N(_0622_),
    .D_N(_0623_),
    .X(_0624_));
 sky130_fd_sc_hd__or4_1 _2352_ (.A(_0614_),
    .B(_0615_),
    .C(_0618_),
    .D(_0624_),
    .X(_0625_));
 sky130_fd_sc_hd__or3_2 _2353_ (.A(\usb2uart.u_usb_cdc.u_sie.crc16_q[7] ),
    .B(_0613_),
    .C(_0625_),
    .X(_0626_));
 sky130_fd_sc_hd__and3_1 _2354_ (.A(_0597_),
    .B(_0588_),
    .C(_0626_),
    .X(_0627_));
 sky130_fd_sc_hd__and4bb_1 _2355_ (.A_N(\usb2uart.u_usb_cdc.u_sie.in_byte_q[1] ),
    .B_N(\usb2uart.u_usb_cdc.u_sie.in_byte_q[0] ),
    .C(_2052_),
    .D(\usb2uart.u_usb_cdc.u_sie.in_byte_q[3] ),
    .X(_0628_));
 sky130_fd_sc_hd__o21a_1 _2356_ (.A1(_2051_),
    .A2(_0628_),
    .B1(_2007_),
    .X(_0629_));
 sky130_fd_sc_hd__inv_2 _2357_ (.A(_0553_),
    .Y(_0630_));
 sky130_fd_sc_hd__a21oi_2 _2358_ (.A1(_2055_),
    .A2(_0629_),
    .B1(_0630_),
    .Y(_0631_));
 sky130_fd_sc_hd__a211o_1 _2359_ (.A1(_0588_),
    .A2(_0596_),
    .B1(_0627_),
    .C1(_0631_),
    .X(_0632_));
 sky130_fd_sc_hd__nand2_2 _2360_ (.A(_2003_),
    .B(_0516_),
    .Y(_0633_));
 sky130_fd_sc_hd__or2_1 _2361_ (.A(\usb2uart.u_usb_cdc.u_sie.phy_state_q[11] ),
    .B(\usb2uart.u_usb_cdc.u_sie.phy_state_q[10] ),
    .X(_0634_));
 sky130_fd_sc_hd__or4_1 _2362_ (.A(_0589_),
    .B(\usb2uart.u_usb_cdc.u_sie.phy_state_q[3] ),
    .C(\usb2uart.u_usb_cdc.u_sie.phy_state_q[2] ),
    .D(\usb2uart.u_usb_cdc.u_sie.phy_state_q[5] ),
    .X(_0635_));
 sky130_fd_sc_hd__o31a_1 _2363_ (.A1(_0528_),
    .A2(_0634_),
    .A3(_0635_),
    .B1(_0516_),
    .X(_0636_));
 sky130_fd_sc_hd__o32a_1 _2364_ (.A1(_0588_),
    .A2(_0633_),
    .A3(_0634_),
    .B1(_0636_),
    .B2(\usb2uart.u_usb_cdc.u_sie.phy_state_q[0] ),
    .X(_0637_));
 sky130_fd_sc_hd__a21o_1 _2365_ (.A1(_0591_),
    .A2(_0632_),
    .B1(_0637_),
    .X(_0017_));
 sky130_fd_sc_hd__or2_1 _2366_ (.A(_2013_),
    .B(_2014_),
    .X(_0638_));
 sky130_fd_sc_hd__clkinv_2 _2367_ (.A(_0453_),
    .Y(_0639_));
 sky130_fd_sc_hd__or2_1 _2368_ (.A(\usb2uart.u_usb_cdc.u_ctrl_endp.byte_cnt_q[0] ),
    .B(\usb2uart.u_usb_cdc.u_ctrl_endp.byte_cnt_q[1] ),
    .X(_0640_));
 sky130_fd_sc_hd__buf_2 _2369_ (.A(_0640_),
    .X(_0641_));
 sky130_fd_sc_hd__or4_1 _2370_ (.A(_0452_),
    .B(_0639_),
    .C(\usb2uart.u_usb_cdc.u_ctrl_endp.req_q[10] ),
    .D(_0641_),
    .X(_0642_));
 sky130_fd_sc_hd__nor2_1 _2371_ (.A(_0455_),
    .B(_0642_),
    .Y(_0643_));
 sky130_fd_sc_hd__and2_2 _2372_ (.A(_2009_),
    .B(_2078_),
    .X(_0644_));
 sky130_fd_sc_hd__inv_2 _2373_ (.A(\usb2uart.u_usb_cdc.u_ctrl_endp.in_req_q ),
    .Y(_0645_));
 sky130_fd_sc_hd__nand2_2 _2374_ (.A(\usb2uart.u_usb_cdc.in_data_ack ),
    .B(_0487_),
    .Y(_0646_));
 sky130_fd_sc_hd__and2b_1 _2375_ (.A_N(_2027_),
    .B(_2043_),
    .X(_0647_));
 sky130_fd_sc_hd__a21o_1 _2376_ (.A1(_0645_),
    .A2(\usb2uart.u_usb_cdc.in_data_ack ),
    .B1(_0647_),
    .X(_0648_));
 sky130_fd_sc_hd__and4_1 _2377_ (.A(_0461_),
    .B(\usb2uart.u_usb_cdc.u_ctrl_endp.state_q[3] ),
    .C(_0487_),
    .D(_0648_),
    .X(_0649_));
 sky130_fd_sc_hd__a31o_1 _2378_ (.A1(_0645_),
    .A2(_2010_),
    .A3(_0646_),
    .B1(_0649_),
    .X(_0650_));
 sky130_fd_sc_hd__a41o_1 _2379_ (.A1(_0497_),
    .A2(_0638_),
    .A3(_0643_),
    .A4(_0644_),
    .B1(_0650_),
    .X(_0651_));
 sky130_fd_sc_hd__a22o_1 _2380_ (.A1(\usb2uart.u_usb_cdc.u_ctrl_endp.state_q[3] ),
    .A2(_0488_),
    .B1(_0651_),
    .B2(_2020_),
    .X(_0016_));
 sky130_fd_sc_hd__clkbuf_4 _2381_ (.A(_2075_),
    .X(_0652_));
 sky130_fd_sc_hd__or3_1 _2382_ (.A(_0652_),
    .B(_0534_),
    .C(_0488_),
    .X(_0653_));
 sky130_fd_sc_hd__inv_2 _2383_ (.A(_0652_),
    .Y(_0654_));
 sky130_fd_sc_hd__nand2_1 _2384_ (.A(_0461_),
    .B(_0647_),
    .Y(_0655_));
 sky130_fd_sc_hd__a22o_1 _2385_ (.A1(_0461_),
    .A2(_2006_),
    .B1(_0655_),
    .B2(\usb2uart.u_usb_cdc.u_ctrl_endp.in_req_q ),
    .X(_0656_));
 sky130_fd_sc_hd__and2b_1 _2386_ (.A_N(_0643_),
    .B(_0497_),
    .X(_0657_));
 sky130_fd_sc_hd__a21o_1 _2387_ (.A1(\usb2uart.u_usb_cdc.u_ctrl_endp.state_q[3] ),
    .A2(_0656_),
    .B1(_0657_),
    .X(_0658_));
 sky130_fd_sc_hd__a31o_1 _2388_ (.A1(_0654_),
    .A2(_0644_),
    .A3(_0658_),
    .B1(\usb2uart.u_usb_cdc.ctrl_stall ),
    .X(_0659_));
 sky130_fd_sc_hd__and2_1 _2389_ (.A(_0653_),
    .B(_0659_),
    .X(_0660_));
 sky130_fd_sc_hd__clkbuf_1 _2390_ (.A(_0660_),
    .X(_0015_));
 sky130_fd_sc_hd__or2_1 _2391_ (.A(_2075_),
    .B(_0487_),
    .X(_0661_));
 sky130_fd_sc_hd__o311a_1 _2392_ (.A1(_0652_),
    .A2(\usb2uart.u_usb_cdc.in_data_ack ),
    .A3(_2017_),
    .B1(_0644_),
    .C1(_0661_),
    .X(_0662_));
 sky130_fd_sc_hd__o21ai_1 _2393_ (.A1(_2012_),
    .A2(_0662_),
    .B1(_0653_),
    .Y(_0014_));
 sky130_fd_sc_hd__a21oi_1 _2394_ (.A1(_0461_),
    .A2(\usb2uart.u_usb_cdc.in_data_ack ),
    .B1(\usb2uart.u_usb_cdc.u_ctrl_endp.in_req_q ),
    .Y(_0663_));
 sky130_fd_sc_hd__o211a_1 _2395_ (.A1(_0461_),
    .A2(\usb2uart.u_usb_cdc.in_data_ack ),
    .B1(_0534_),
    .C1(_0663_),
    .X(_0664_));
 sky130_fd_sc_hd__a31o_1 _2396_ (.A1(_0487_),
    .A2(_0655_),
    .A3(_0664_),
    .B1(_0652_),
    .X(_0665_));
 sky130_fd_sc_hd__nor2_1 _2397_ (.A(_2017_),
    .B(_0646_),
    .Y(_0666_));
 sky130_fd_sc_hd__a22o_1 _2398_ (.A1(_0652_),
    .A2(_0473_),
    .B1(_2082_),
    .B2(_0666_),
    .X(_0667_));
 sky130_fd_sc_hd__a21oi_1 _2399_ (.A1(\usb2uart.u_usb_cdc.u_ctrl_endp.state_q[3] ),
    .A2(_0665_),
    .B1(_0667_),
    .Y(_0668_));
 sky130_fd_sc_hd__a2bb2o_1 _2400_ (.A1_N(_0668_),
    .A2_N(_0488_),
    .B1(\usb2uart.u_usb_cdc.u_ctrl_endp.state_q[0] ),
    .B2(_0653_),
    .X(_0013_));
 sky130_fd_sc_hd__inv_2 _2401_ (.A(_0507_),
    .Y(_0669_));
 sky130_fd_sc_hd__or3b_1 _2402_ (.A(_0468_),
    .B(\usb2uart.u_usb_cdc.out_data[0] ),
    .C_N(\usb2uart.u_usb_cdc.out_data[1] ),
    .X(_0670_));
 sky130_fd_sc_hd__or2_1 _2403_ (.A(_0483_),
    .B(_0670_),
    .X(_0671_));
 sky130_fd_sc_hd__inv_2 _2404_ (.A(_0671_),
    .Y(_0672_));
 sky130_fd_sc_hd__inv_2 _2405_ (.A(\usb2uart.u_usb_cdc.u_ctrl_endp.dev_state_qq[0] ),
    .Y(_0673_));
 sky130_fd_sc_hd__o21ai_1 _2406_ (.A1(_0673_),
    .A2(\usb2uart.u_usb_cdc.u_ctrl_endp.dev_state_qq[1] ),
    .B1(\usb2uart.u_usb_cdc.u_ctrl_endp.in_dir_q ),
    .Y(_0674_));
 sky130_fd_sc_hd__and3b_1 _2407_ (.A_N(_0674_),
    .B(_2002_),
    .C(_0485_),
    .X(_0675_));
 sky130_fd_sc_hd__a32o_1 _2408_ (.A1(\usb2uart.u_usb_cdc.u_ctrl_endp.req_q[11] ),
    .A2(_0669_),
    .A3(_0672_),
    .B1(_0675_),
    .B2(_0459_),
    .X(_0676_));
 sky130_fd_sc_hd__or2b_1 _2409_ (.A(\usb2uart.u_usb_cdc.u_ctrl_endp.rec_q[0] ),
    .B_N(\usb2uart.u_usb_cdc.u_ctrl_endp.rec_q[1] ),
    .X(_0677_));
 sky130_fd_sc_hd__clkinv_2 _2410_ (.A(\usb2uart.u_usb_cdc.out_data[7] ),
    .Y(_0678_));
 sky130_fd_sc_hd__o21a_1 _2411_ (.A1(_0482_),
    .A2(_0678_),
    .B1(_0465_),
    .X(_0679_));
 sky130_fd_sc_hd__or4_2 _2412_ (.A(_0483_),
    .B(_0467_),
    .C(_0677_),
    .D(_0679_),
    .X(_0680_));
 sky130_fd_sc_hd__nor3_4 _2413_ (.A(_0465_),
    .B(_0483_),
    .C(_0468_),
    .Y(_0681_));
 sky130_fd_sc_hd__or3b_1 _2414_ (.A(\usb2uart.u_usb_cdc.out_data[4] ),
    .B(\usb2uart.u_usb_cdc.u_ctrl_endp.rec_q[1] ),
    .C_N(\usb2uart.u_usb_cdc.u_ctrl_endp.rec_q[0] ),
    .X(_0682_));
 sky130_fd_sc_hd__o21ai_1 _2415_ (.A1(_0482_),
    .A2(_0462_),
    .B1(_0682_),
    .Y(_0683_));
 sky130_fd_sc_hd__nand2_1 _2416_ (.A(_0681_),
    .B(_0683_),
    .Y(_0684_));
 sky130_fd_sc_hd__nand2_1 _2417_ (.A(_0680_),
    .B(_0684_),
    .Y(_0685_));
 sky130_fd_sc_hd__and3_1 _2418_ (.A(_0473_),
    .B(_0495_),
    .C(_0685_),
    .X(_0686_));
 sky130_fd_sc_hd__and3_1 _2419_ (.A(_2009_),
    .B(_2020_),
    .C(_2078_),
    .X(_0687_));
 sky130_fd_sc_hd__nor2_4 _2420_ (.A(_2012_),
    .B(_0487_),
    .Y(_0688_));
 sky130_fd_sc_hd__and3_1 _2421_ (.A(_0456_),
    .B(_0687_),
    .C(_0688_),
    .X(_0689_));
 sky130_fd_sc_hd__or3b_4 _2422_ (.A(_0498_),
    .B(_0497_),
    .C_N(_0687_),
    .X(_0690_));
 sky130_fd_sc_hd__and3_1 _2423_ (.A(_2079_),
    .B(_0485_),
    .C(_0479_),
    .X(_0691_));
 sky130_fd_sc_hd__nor2_1 _2424_ (.A(_0474_),
    .B(_0489_),
    .Y(_0692_));
 sky130_fd_sc_hd__or2_1 _2425_ (.A(_0481_),
    .B(_0504_),
    .X(_0693_));
 sky130_fd_sc_hd__o211a_1 _2426_ (.A1(_0692_),
    .A2(_0693_),
    .B1(_2079_),
    .C1(_0485_),
    .X(_0694_));
 sky130_fd_sc_hd__or4_2 _2427_ (.A(_0689_),
    .B(_0690_),
    .C(_0691_),
    .D(_0694_),
    .X(_0695_));
 sky130_fd_sc_hd__o21a_1 _2428_ (.A1(_0686_),
    .A2(_0695_),
    .B1(\usb2uart.u_usb_cdc.u_ctrl_endp.req_q[11] ),
    .X(_0696_));
 sky130_fd_sc_hd__a21o_1 _2429_ (.A1(_2080_),
    .A2(_0676_),
    .B1(_0696_),
    .X(_0003_));
 sky130_fd_sc_hd__or2_1 _2430_ (.A(_0456_),
    .B(_0493_),
    .X(_0697_));
 sky130_fd_sc_hd__a31o_1 _2431_ (.A1(_0687_),
    .A2(_0688_),
    .A3(_0697_),
    .B1(_0690_),
    .X(_0698_));
 sky130_fd_sc_hd__nand2_2 _2432_ (.A(_0464_),
    .B(_0681_),
    .Y(_0699_));
 sky130_fd_sc_hd__buf_2 _2433_ (.A(\usb2uart.u_usb_cdc.u_ctrl_endp.req_q[8] ),
    .X(_0700_));
 sky130_fd_sc_hd__or2_1 _2434_ (.A(\usb2uart.u_usb_cdc.u_ctrl_endp.req_q[2] ),
    .B(_0700_),
    .X(_0701_));
 sky130_fd_sc_hd__nor2_1 _2435_ (.A(\usb2uart.u_usb_cdc.u_ctrl_endp.req_q[1] ),
    .B(\usb2uart.u_usb_cdc.u_ctrl_endp.req_q[7] ),
    .Y(_0702_));
 sky130_fd_sc_hd__or3b_1 _2436_ (.A(\usb2uart.u_usb_cdc.u_ctrl_endp.req_q[3] ),
    .B(_0701_),
    .C_N(_0702_),
    .X(_0703_));
 sky130_fd_sc_hd__a22o_1 _2437_ (.A1(\usb2uart.u_usb_cdc.u_ctrl_endp.req_q[5] ),
    .A2(_0484_),
    .B1(_0699_),
    .B2(_0703_),
    .X(_0704_));
 sky130_fd_sc_hd__and3_1 _2438_ (.A(\usb2uart.u_usb_cdc.u_ctrl_endp.req_q[11] ),
    .B(_0680_),
    .C(_0684_),
    .X(_0705_));
 sky130_fd_sc_hd__a211o_1 _2439_ (.A1(\usb2uart.u_usb_cdc.u_ctrl_endp.req_q[6] ),
    .A2(_0680_),
    .B1(_0704_),
    .C1(_0705_),
    .X(_0706_));
 sky130_fd_sc_hd__a2111o_1 _2440_ (.A1(_0482_),
    .A2(_0465_),
    .B1(\usb2uart.u_usb_cdc.out_data[4] ),
    .C1(_0466_),
    .D1(_0483_),
    .X(_0707_));
 sky130_fd_sc_hd__and4_1 _2441_ (.A(_0473_),
    .B(_0492_),
    .C(_0457_),
    .D(_0707_),
    .X(_0708_));
 sky130_fd_sc_hd__and2_2 _2442_ (.A(\usb2uart.u_usb_cdc.u_ctrl_endp.dev_state_qq[0] ),
    .B(\usb2uart.u_usb_cdc.u_ctrl_endp.dev_state_qq[1] ),
    .X(_0709_));
 sky130_fd_sc_hd__and4b_1 _2443_ (.A_N(_0466_),
    .B(_0678_),
    .C(\usb2uart.u_usb_cdc.u_ctrl_endp.class_q ),
    .D(\usb2uart.u_usb_cdc.out_data[5] ),
    .X(_0710_));
 sky130_fd_sc_hd__and4bb_1 _2444_ (.A_N(\usb2uart.u_usb_cdc.out_data[4] ),
    .B_N(_0483_),
    .C(_0709_),
    .D(_0710_),
    .X(_0711_));
 sky130_fd_sc_hd__o21ba_1 _2445_ (.A1(_0673_),
    .A2(\usb2uart.u_usb_cdc.u_ctrl_endp.dev_state_qq[1] ),
    .B1_N(\usb2uart.u_usb_cdc.u_ctrl_endp.in_dir_q ),
    .X(_0712_));
 sky130_fd_sc_hd__nand2_1 _2446_ (.A(_0482_),
    .B(_0681_),
    .Y(_0713_));
 sky130_fd_sc_hd__or3_1 _2447_ (.A(\usb2uart.u_usb_cdc.out_data[2] ),
    .B(_0469_),
    .C(_0468_),
    .X(_0714_));
 sky130_fd_sc_hd__or3_1 _2448_ (.A(_0464_),
    .B(_0465_),
    .C(_0714_),
    .X(_0715_));
 sky130_fd_sc_hd__or3b_1 _2449_ (.A(\usb2uart.u_usb_cdc.u_ctrl_endp.class_q ),
    .B(_0462_),
    .C_N(_0712_),
    .X(_0716_));
 sky130_fd_sc_hd__a21bo_1 _2450_ (.A1(_2002_),
    .A2(_0715_),
    .B1_N(_0716_),
    .X(_0717_));
 sky130_fd_sc_hd__and4b_1 _2451_ (.A_N(\usb2uart.u_usb_cdc.u_ctrl_endp.rec_q[1] ),
    .B(_0709_),
    .C(_0461_),
    .D(\usb2uart.u_usb_cdc.u_ctrl_endp.rec_q[0] ),
    .X(_0718_));
 sky130_fd_sc_hd__or3_1 _2452_ (.A(\usb2uart.u_usb_cdc.out_data[2] ),
    .B(_0469_),
    .C(_0670_),
    .X(_0719_));
 sky130_fd_sc_hd__nand2_1 _2453_ (.A(_0485_),
    .B(_0674_),
    .Y(_0720_));
 sky130_fd_sc_hd__o221a_1 _2454_ (.A1(_0463_),
    .A2(_0471_),
    .B1(_0718_),
    .B2(_0719_),
    .C1(_0720_),
    .X(_0721_));
 sky130_fd_sc_hd__o211a_1 _2455_ (.A1(_0712_),
    .A2(_0713_),
    .B1(_0717_),
    .C1(_0721_),
    .X(_0722_));
 sky130_fd_sc_hd__nor2_1 _2456_ (.A(_0711_),
    .B(_0722_),
    .Y(_0723_));
 sky130_fd_sc_hd__or3_1 _2457_ (.A(\usb2uart.u_usb_cdc.u_ctrl_endp.req_q[5] ),
    .B(\usb2uart.u_usb_cdc.u_ctrl_endp.req_q[11] ),
    .C(\usb2uart.u_usb_cdc.u_ctrl_endp.req_q[6] ),
    .X(_0724_));
 sky130_fd_sc_hd__or2_1 _2458_ (.A(\usb2uart.u_usb_cdc.u_ctrl_endp.req_q[9] ),
    .B(_0724_),
    .X(_0725_));
 sky130_fd_sc_hd__or4_1 _2459_ (.A(\usb2uart.u_usb_cdc.u_ctrl_endp.req_q[10] ),
    .B(\usb2uart.u_usb_cdc.u_ctrl_endp.req_q[4] ),
    .C(_0725_),
    .D(_0703_),
    .X(_0726_));
 sky130_fd_sc_hd__nor2_1 _2460_ (.A(\usb2uart.u_usb_cdc.u_ctrl_endp.rec_q[0] ),
    .B(\usb2uart.u_usb_cdc.u_ctrl_endp.rec_q[1] ),
    .Y(_0727_));
 sky130_fd_sc_hd__nor2_1 _2461_ (.A(_0470_),
    .B(_0670_),
    .Y(_0728_));
 sky130_fd_sc_hd__a31o_1 _2462_ (.A1(_0461_),
    .A2(_0727_),
    .A3(_0728_),
    .B1(\usb2uart.u_usb_cdc.u_ctrl_endp.class_q ),
    .X(_0729_));
 sky130_fd_sc_hd__or4_1 _2463_ (.A(\usb2uart.u_usb_cdc.out_data[0] ),
    .B(_0465_),
    .C(_0462_),
    .D(_0674_),
    .X(_0730_));
 sky130_fd_sc_hd__o211a_1 _2464_ (.A1(_0714_),
    .A2(_0730_),
    .B1(_0715_),
    .C1(_0719_),
    .X(_0731_));
 sky130_fd_sc_hd__and4b_1 _2465_ (.A_N(_0729_),
    .B(_0471_),
    .C(_0484_),
    .D(_0731_),
    .X(_0732_));
 sky130_fd_sc_hd__o311a_1 _2466_ (.A1(_0723_),
    .A2(_0726_),
    .A3(_0732_),
    .B1(_0458_),
    .C1(_0473_),
    .X(_0733_));
 sky130_fd_sc_hd__a311o_1 _2467_ (.A1(_0473_),
    .A2(_0495_),
    .A3(_0706_),
    .B1(_0708_),
    .C1(_0733_),
    .X(_0734_));
 sky130_fd_sc_hd__inv_2 _2468_ (.A(\usb2uart.u_usb_cdc.u_ctrl_endp.req_q[1] ),
    .Y(_0735_));
 sky130_fd_sc_hd__nor2_1 _2469_ (.A(\usb2uart.u_usb_cdc.u_ctrl_endp.req_q[7] ),
    .B(\usb2uart.u_usb_cdc.u_ctrl_endp.req_q[6] ),
    .Y(_0736_));
 sky130_fd_sc_hd__nand2_1 _2470_ (.A(_0735_),
    .B(_0736_),
    .Y(_0737_));
 sky130_fd_sc_hd__or3b_1 _2471_ (.A(\usb2uart.u_usb_cdc.u_ctrl_endp.req_q[3] ),
    .B(_0724_),
    .C_N(_0702_),
    .X(_0738_));
 sky130_fd_sc_hd__a22o_1 _2472_ (.A1(_0508_),
    .A2(_0737_),
    .B1(_0738_),
    .B2(_0693_),
    .X(_0739_));
 sky130_fd_sc_hd__or3_1 _2473_ (.A(_0504_),
    .B(_0669_),
    .C(_0692_),
    .X(_0740_));
 sky130_fd_sc_hd__a31o_1 _2474_ (.A1(\usb2uart.u_usb_cdc.u_ctrl_endp.req_q[9] ),
    .A2(_0671_),
    .A3(_0713_),
    .B1(\usb2uart.u_usb_cdc.u_ctrl_endp.req_q[10] ),
    .X(_0741_));
 sky130_fd_sc_hd__a22o_1 _2475_ (.A1(\usb2uart.u_usb_cdc.u_ctrl_endp.req_q[10] ),
    .A2(_0740_),
    .B1(_0741_),
    .B2(_0481_),
    .X(_0742_));
 sky130_fd_sc_hd__or2_1 _2476_ (.A(\usb2uart.u_usb_cdc.u_ctrl_endp.req_q[3] ),
    .B(_0725_),
    .X(_0743_));
 sky130_fd_sc_hd__a22o_1 _2477_ (.A1(\usb2uart.u_usb_cdc.u_ctrl_endp.req_q[7] ),
    .A2(_0484_),
    .B1(_0699_),
    .B2(_0743_),
    .X(_0744_));
 sky130_fd_sc_hd__a221o_1 _2478_ (.A1(\usb2uart.u_usb_cdc.out_data[7] ),
    .A2(\usb2uart.u_usb_cdc.u_ctrl_endp.req_q[1] ),
    .B1(\usb2uart.u_usb_cdc.u_ctrl_endp.req_q[6] ),
    .B2(_0677_),
    .C1(_0744_),
    .X(_0745_));
 sky130_fd_sc_hd__a22o_1 _2479_ (.A1(\usb2uart.u_usb_cdc.u_ctrl_endp.req_q[11] ),
    .A2(_0671_),
    .B1(_0713_),
    .B2(_0505_),
    .X(_0746_));
 sky130_fd_sc_hd__o41a_1 _2480_ (.A1(\usb2uart.u_usb_cdc.u_ctrl_endp.req_q[11] ),
    .A2(_0505_),
    .A3(_0701_),
    .A4(_0737_),
    .B1(_0699_),
    .X(_0747_));
 sky130_fd_sc_hd__o21a_1 _2481_ (.A1(\usb2uart.u_usb_cdc.u_ctrl_endp.req_q[10] ),
    .A2(_0747_),
    .B1(_0479_),
    .X(_0748_));
 sky130_fd_sc_hd__a221o_1 _2482_ (.A1(_0692_),
    .A2(_0745_),
    .B1(_0746_),
    .B2(_0669_),
    .C1(_0748_),
    .X(_0749_));
 sky130_fd_sc_hd__a211o_1 _2483_ (.A1(_0699_),
    .A2(_0739_),
    .B1(_0742_),
    .C1(_0749_),
    .X(_0750_));
 sky130_fd_sc_hd__a21o_1 _2484_ (.A1(_2020_),
    .A2(_0734_),
    .B1(_0750_),
    .X(_0751_));
 sky130_fd_sc_hd__a22o_1 _2485_ (.A1(\usb2uart.u_usb_cdc.u_ctrl_endp.req_q[10] ),
    .A2(_0698_),
    .B1(_0751_),
    .B2(_2080_),
    .X(_0002_));
 sky130_fd_sc_hd__and3_1 _2486_ (.A(_2080_),
    .B(_0485_),
    .C(_0692_),
    .X(_0752_));
 sky130_fd_sc_hd__o31a_1 _2487_ (.A1(_0479_),
    .A2(_0504_),
    .A3(_0669_),
    .B1(_2080_),
    .X(_0753_));
 sky130_fd_sc_hd__o31a_1 _2488_ (.A1(_0752_),
    .A2(_0698_),
    .A3(_0753_),
    .B1(\usb2uart.u_usb_cdc.u_ctrl_endp.req_q[9] ),
    .X(_0754_));
 sky130_fd_sc_hd__a41o_1 _2489_ (.A1(_0461_),
    .A2(_0460_),
    .A3(_0727_),
    .A4(_0728_),
    .B1(_0754_),
    .X(_0012_));
 sky130_fd_sc_hd__nand2_1 _2490_ (.A(_2080_),
    .B(_0481_),
    .Y(_0755_));
 sky130_fd_sc_hd__or4bb_1 _2491_ (.A(_0496_),
    .B(_0500_),
    .C_N(_0755_),
    .D_N(_0490_),
    .X(_0756_));
 sky130_fd_sc_hd__nor2_1 _2492_ (.A(_0477_),
    .B(_0476_),
    .Y(_0757_));
 sky130_fd_sc_hd__a211o_1 _2493_ (.A1(_0757_),
    .A2(_0688_),
    .B1(_0511_),
    .C1(_0691_),
    .X(_0758_));
 sky130_fd_sc_hd__inv_2 _2494_ (.A(_0755_),
    .Y(_0759_));
 sky130_fd_sc_hd__clkbuf_4 _2495_ (.A(_0700_),
    .X(_0760_));
 sky130_fd_sc_hd__a31o_1 _2496_ (.A1(\usb2uart.u_usb_cdc.u_ctrl_endp.req_q[9] ),
    .A2(_0759_),
    .A3(_0672_),
    .B1(_0760_),
    .X(_0761_));
 sky130_fd_sc_hd__o21a_1 _2497_ (.A1(_0756_),
    .A2(_0758_),
    .B1(_0761_),
    .X(_0011_));
 sky130_fd_sc_hd__and3_1 _2498_ (.A(\usb2uart.u_usb_cdc.u_ctrl_endp.req_q[0] ),
    .B(_0688_),
    .C(_0458_),
    .X(_0762_));
 sky130_fd_sc_hd__nor2_1 _2499_ (.A(_0716_),
    .B(_0715_),
    .Y(_0763_));
 sky130_fd_sc_hd__a21oi_1 _2500_ (.A1(_0490_),
    .A2(_0755_),
    .B1(_0699_),
    .Y(_0764_));
 sky130_fd_sc_hd__or2_1 _2501_ (.A(_0511_),
    .B(_0691_),
    .X(_0765_));
 sky130_fd_sc_hd__or4_1 _2502_ (.A(_0464_),
    .B(_0465_),
    .C(_0483_),
    .D(_0468_),
    .X(_0766_));
 sky130_fd_sc_hd__nor2_1 _2503_ (.A(_0490_),
    .B(_0766_),
    .Y(_0767_));
 sky130_fd_sc_hd__o41a_1 _2504_ (.A1(_0510_),
    .A2(_0764_),
    .A3(_0765_),
    .A4(_0767_),
    .B1(\usb2uart.u_usb_cdc.u_ctrl_endp.req_q[7] ),
    .X(_0768_));
 sky130_fd_sc_hd__a31o_1 _2505_ (.A1(_0687_),
    .A2(_0762_),
    .A3(_0763_),
    .B1(_0768_),
    .X(_0010_));
 sky130_fd_sc_hd__nor2_1 _2506_ (.A(_0464_),
    .B(_0484_),
    .Y(_0769_));
 sky130_fd_sc_hd__nor3_1 _2507_ (.A(_0699_),
    .B(_0490_),
    .C(_0677_),
    .Y(_0770_));
 sky130_fd_sc_hd__or2_1 _2508_ (.A(_0500_),
    .B(_0509_),
    .X(_0771_));
 sky130_fd_sc_hd__and3_1 _2509_ (.A(_2079_),
    .B(_0485_),
    .C(_0481_),
    .X(_0772_));
 sky130_fd_sc_hd__nand2_1 _2510_ (.A(_2006_),
    .B(_0495_),
    .Y(_0773_));
 sky130_fd_sc_hd__or3_1 _2511_ (.A(_0474_),
    .B(_0773_),
    .C(_0680_),
    .X(_0774_));
 sky130_fd_sc_hd__or4b_1 _2512_ (.A(_0511_),
    .B(_0691_),
    .C(_0772_),
    .D_N(_0774_),
    .X(_0775_));
 sky130_fd_sc_hd__o31a_1 _2513_ (.A1(_0770_),
    .A2(_0771_),
    .A3(_0775_),
    .B1(\usb2uart.u_usb_cdc.u_ctrl_endp.req_q[6] ),
    .X(_0776_));
 sky130_fd_sc_hd__a31o_1 _2514_ (.A1(_0460_),
    .A2(_0712_),
    .A3(_0769_),
    .B1(_0776_),
    .X(_0009_));
 sky130_fd_sc_hd__nor2_1 _2515_ (.A(\usb2uart.u_usb_cdc.u_sie.phy_state_q[7] ),
    .B(_0553_),
    .Y(_0777_));
 sky130_fd_sc_hd__nor2_1 _2516_ (.A(\usb2uart.u_usb_cdc.u_sie.rx_err ),
    .B(_0777_),
    .Y(_0778_));
 sky130_fd_sc_hd__nand2_1 _2517_ (.A(_2049_),
    .B(_0778_),
    .Y(_0779_));
 sky130_fd_sc_hd__inv_2 _2518_ (.A(_0779_),
    .Y(\usb2uart.u_usb_cdc.bulk_in_req ));
 sky130_fd_sc_hd__clkbuf_4 _2519_ (.A(_2061_),
    .X(_0780_));
 sky130_fd_sc_hd__buf_2 _2520_ (.A(\usb2uart.u_usb_cdc.u_sie.u_phy_tx.tx_valid_q ),
    .X(_0781_));
 sky130_fd_sc_hd__nor2_2 _2521_ (.A(_0781_),
    .B(_2063_),
    .Y(_0782_));
 sky130_fd_sc_hd__nand2_2 _2522_ (.A(\usb2uart.u_usb_cdc.u_sie.u_phy_tx.clk_cnt_q[1] ),
    .B(\usb2uart.u_usb_cdc.u_sie.u_phy_tx.clk_cnt_q[0] ),
    .Y(_0783_));
 sky130_fd_sc_hd__nand2b_1 _2523_ (.A_N(_0783_),
    .B(_2060_),
    .Y(_0784_));
 sky130_fd_sc_hd__buf_2 _2524_ (.A(_2063_),
    .X(_0785_));
 sky130_fd_sc_hd__or2_1 _2525_ (.A(_0784_),
    .B(_0785_),
    .X(_0786_));
 sky130_fd_sc_hd__a32o_1 _2526_ (.A1(\usb2uart.u_usb_cdc.u_sie.u_phy_tx.tx_state_q[1] ),
    .A2(_0780_),
    .A3(_0782_),
    .B1(_0786_),
    .B2(\usb2uart.u_usb_cdc.u_sie.u_phy_tx.tx_state_q[3] ),
    .X(_0037_));
 sky130_fd_sc_hd__inv_2 _2527_ (.A(net6),
    .Y(_0787_));
 sky130_fd_sc_hd__a2bb2o_1 _2528_ (.A1_N(_0787_),
    .A2_N(_2062_),
    .B1(_0786_),
    .B2(\usb2uart.u_usb_cdc.u_sie.u_phy_tx.tx_state_q[2] ),
    .X(_0036_));
 sky130_fd_sc_hd__buf_2 _2529_ (.A(_0784_),
    .X(_0788_));
 sky130_fd_sc_hd__nor2_1 _2530_ (.A(_0788_),
    .B(_0785_),
    .Y(_0789_));
 sky130_fd_sc_hd__or2_1 _2531_ (.A(\usb2uart.u_usb_cdc.u_sie.u_phy_tx.tx_valid_q ),
    .B(_2063_),
    .X(_0790_));
 sky130_fd_sc_hd__or2_1 _2532_ (.A(\usb2uart.u_usb_cdc.u_sie.u_phy_tx.tx_state_q[1] ),
    .B(\usb2uart.u_usb_cdc.u_sie.u_phy_tx.tx_state_q[2] ),
    .X(_0791_));
 sky130_fd_sc_hd__o221a_1 _2533_ (.A1(\usb2uart.u_usb_cdc.u_sie.u_phy_tx.tx_state_q[1] ),
    .A2(_0789_),
    .B1(_0790_),
    .B2(_0788_),
    .C1(_0791_),
    .X(_0035_));
 sky130_fd_sc_hd__inv_2 _2534_ (.A(\usb2uart.u_usb_cdc.u_sie.u_phy_tx.tx_state_q[3] ),
    .Y(_0792_));
 sky130_fd_sc_hd__nand2_1 _2535_ (.A(_0781_),
    .B(_0792_),
    .Y(_0793_));
 sky130_fd_sc_hd__or2_1 _2536_ (.A(\usb2uart.u_usb_cdc.u_sie.u_phy_tx.tx_state_q[3] ),
    .B(\usb2uart.u_usb_cdc.u_sie.u_phy_tx.tx_state_q[2] ),
    .X(_0794_));
 sky130_fd_sc_hd__a32o_1 _2537_ (.A1(_0789_),
    .A2(_0793_),
    .A3(_0794_),
    .B1(_2062_),
    .B2(net6),
    .X(_0034_));
 sky130_fd_sc_hd__clkbuf_4 _2538_ (.A(_2070_),
    .X(_0795_));
 sky130_fd_sc_hd__o311ai_4 _2539_ (.A1(\usb2uart.u_usb_cdc.u_ctrl_endp.dev_state_qq[0] ),
    .A2(\usb2uart.u_usb_cdc.u_ctrl_endp.dev_state_qq[1] ),
    .A3(\usb2uart.u_usb_cdc.u_ctrl_endp.usb_reset_q ),
    .B1(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.rx_en_q ),
    .C1(net6),
    .Y(_0796_));
 sky130_fd_sc_hd__nor2_1 _2540_ (.A(_0795_),
    .B(_0796_),
    .Y(_0797_));
 sky130_fd_sc_hd__or4_1 _2541_ (.A(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.data_q[0] ),
    .B(\usb2uart.u_usb_cdc.u_sie.rx_data[0] ),
    .C(\usb2uart.u_usb_cdc.u_sie.rx_data[1] ),
    .D(\usb2uart.u_usb_cdc.u_sie.rx_data[3] ),
    .X(_0798_));
 sky130_fd_sc_hd__or2_4 _2542_ (.A(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.nrzi_q[2] ),
    .B(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.nrzi_q[3] ),
    .X(_0799_));
 sky130_fd_sc_hd__nor4_1 _2543_ (.A(\usb2uart.u_usb_cdc.u_sie.rx_data[2] ),
    .B(\usb2uart.u_usb_cdc.u_sie.rx_data[4] ),
    .C(_0798_),
    .D(_0799_),
    .Y(_0800_));
 sky130_fd_sc_hd__and4b_1 _2544_ (.A_N(\usb2uart.u_usb_cdc.u_sie.rx_data[5] ),
    .B(\usb2uart.u_usb_cdc.u_sie.rx_data[6] ),
    .C(\usb2uart.u_usb_cdc.u_sie.rx_data[7] ),
    .D(_0800_),
    .X(_0801_));
 sky130_fd_sc_hd__and2_1 _2545_ (.A(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.rx_state_q[4] ),
    .B(_0795_),
    .X(_0802_));
 sky130_fd_sc_hd__a31o_1 _2546_ (.A1(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.rx_state_q[2] ),
    .A2(_0797_),
    .A3(_0801_),
    .B1(_0802_),
    .X(_0033_));
 sky130_fd_sc_hd__nand2_1 _2547_ (.A(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.nrzi_q[2] ),
    .B(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.nrzi_q[3] ),
    .Y(_0803_));
 sky130_fd_sc_hd__and2_1 _2548_ (.A(_0799_),
    .B(_0803_),
    .X(_0804_));
 sky130_fd_sc_hd__or2_1 _2549_ (.A(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.nrzi_q[3] ),
    .B(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.nrzi_q[1] ),
    .X(_0805_));
 sky130_fd_sc_hd__nand2_1 _2550_ (.A(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.nrzi_q[3] ),
    .B(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.nrzi_q[1] ),
    .Y(_0806_));
 sky130_fd_sc_hd__and2b_1 _2551_ (.A_N(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.nrzi_q[2] ),
    .B(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.nrzi_q[0] ),
    .X(_0807_));
 sky130_fd_sc_hd__and2b_1 _2552_ (.A_N(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.nrzi_q[0] ),
    .B(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.nrzi_q[2] ),
    .X(_0808_));
 sky130_fd_sc_hd__a211o_1 _2553_ (.A1(_0805_),
    .A2(_0806_),
    .B1(_0807_),
    .C1(_0808_),
    .X(_0809_));
 sky130_fd_sc_hd__and2_1 _2554_ (.A(_0804_),
    .B(_0809_),
    .X(_0810_));
 sky130_fd_sc_hd__or4b_1 _2555_ (.A(_2067_),
    .B(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.nrzi_q[1] ),
    .C(_2070_),
    .D_N(_0807_),
    .X(_0811_));
 sky130_fd_sc_hd__nor2_1 _2556_ (.A(_0796_),
    .B(_0811_),
    .Y(_0812_));
 sky130_fd_sc_hd__a22o_1 _2557_ (.A1(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.rx_state_q[3] ),
    .A2(_0795_),
    .B1(_0812_),
    .B2(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.rx_state_q[0] ),
    .X(_0813_));
 sky130_fd_sc_hd__a31o_1 _2558_ (.A1(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.rx_state_q[3] ),
    .A2(_0797_),
    .A3(_0810_),
    .B1(_0813_),
    .X(_0032_));
 sky130_fd_sc_hd__or4_1 _2559_ (.A(\usb2uart.u_usb_cdc.u_sie.rx_data[3] ),
    .B(\usb2uart.u_usb_cdc.u_sie.rx_data[5] ),
    .C(\usb2uart.u_usb_cdc.u_sie.rx_data[6] ),
    .D(\usb2uart.u_usb_cdc.u_sie.rx_data[7] ),
    .X(_0814_));
 sky130_fd_sc_hd__or4_1 _2560_ (.A(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.nrzi_q[2] ),
    .B(_2067_),
    .C(\usb2uart.u_usb_cdc.u_sie.rx_data[2] ),
    .D(\usb2uart.u_usb_cdc.u_sie.rx_data[4] ),
    .X(_0815_));
 sky130_fd_sc_hd__nor2_1 _2561_ (.A(_0814_),
    .B(_0815_),
    .Y(_0816_));
 sky130_fd_sc_hd__nand2_1 _2562_ (.A(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.rx_state_q[3] ),
    .B(_0816_),
    .Y(_0817_));
 sky130_fd_sc_hd__nor2_1 _2563_ (.A(_0809_),
    .B(_0817_),
    .Y(_0818_));
 sky130_fd_sc_hd__nand2_1 _2564_ (.A(_0804_),
    .B(_0809_),
    .Y(_0819_));
 sky130_fd_sc_hd__nor2_1 _2565_ (.A(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.nrzi_q[1] ),
    .B(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.nrzi_q[0] ),
    .Y(_0820_));
 sky130_fd_sc_hd__or2_1 _2566_ (.A(_2065_),
    .B(_0820_),
    .X(_0821_));
 sky130_fd_sc_hd__clkinv_2 _2567_ (.A(_0821_),
    .Y(_0822_));
 sky130_fd_sc_hd__a2bb2o_1 _2568_ (.A1_N(_2066_),
    .A2_N(_0799_),
    .B1(_0804_),
    .B2(_0822_),
    .X(_0823_));
 sky130_fd_sc_hd__o21ba_1 _2569_ (.A1(_0819_),
    .A2(_0820_),
    .B1_N(_0823_),
    .X(_0824_));
 sky130_fd_sc_hd__and2b_1 _2570_ (.A_N(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.clk_cnt_q[1] ),
    .B(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.clk_cnt_q[0] ),
    .X(_0825_));
 sky130_fd_sc_hd__clkbuf_4 _2571_ (.A(_0825_),
    .X(_0826_));
 sky130_fd_sc_hd__o21ai_1 _2572_ (.A1(_0796_),
    .A2(_0824_),
    .B1(_0826_),
    .Y(_0827_));
 sky130_fd_sc_hd__nand2_1 _2573_ (.A(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.rx_state_q[2] ),
    .B(_0827_),
    .Y(_0828_));
 sky130_fd_sc_hd__a21bo_1 _2574_ (.A1(_0797_),
    .A2(_0818_),
    .B1_N(_0828_),
    .X(_0031_));
 sky130_fd_sc_hd__inv_2 _2575_ (.A(_0801_),
    .Y(_0829_));
 sky130_fd_sc_hd__nand2_1 _2576_ (.A(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.nrzi_q[2] ),
    .B(_2067_),
    .Y(_0830_));
 sky130_fd_sc_hd__a32o_1 _2577_ (.A1(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.rx_state_q[2] ),
    .A2(_0829_),
    .A3(_0824_),
    .B1(_0830_),
    .B2(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.rx_state_q[4] ),
    .X(_0831_));
 sky130_fd_sc_hd__a22o_1 _2578_ (.A1(_0589_),
    .A2(_0795_),
    .B1(_0797_),
    .B2(_0831_),
    .X(_0030_));
 sky130_fd_sc_hd__nand2_1 _2579_ (.A(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.rx_state_q[3] ),
    .B(_0819_),
    .Y(_0832_));
 sky130_fd_sc_hd__nor2_1 _2580_ (.A(_0816_),
    .B(_0832_),
    .Y(_0833_));
 sky130_fd_sc_hd__or3_1 _2581_ (.A(_2068_),
    .B(_0796_),
    .C(_0833_),
    .X(_0834_));
 sky130_fd_sc_hd__a22o_1 _2582_ (.A1(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.rx_state_q[0] ),
    .A2(_0811_),
    .B1(_0834_),
    .B2(_0826_),
    .X(_0029_));
 sky130_fd_sc_hd__inv_2 _2583_ (.A(\usb2uart.u_usb_cdc.u_sie.phy_state_q[11] ),
    .Y(_0835_));
 sky130_fd_sc_hd__buf_2 _2584_ (.A(_0516_),
    .X(_0836_));
 sky130_fd_sc_hd__nand2_1 _2585_ (.A(_0597_),
    .B(_0588_),
    .Y(_0837_));
 sky130_fd_sc_hd__or3_2 _2586_ (.A(_0633_),
    .B(_0837_),
    .C(_0626_),
    .X(_0838_));
 sky130_fd_sc_hd__o21ai_1 _2587_ (.A1(_0835_),
    .A2(_0836_),
    .B1(_0838_),
    .Y(_0019_));
 sky130_fd_sc_hd__a22o_1 _2588_ (.A1(\usb2uart.u_usb_cdc.u_sie.phy_state_q[10] ),
    .A2(_0515_),
    .B1(_0591_),
    .B2(\usb2uart.u_usb_cdc.u_sie.phy_state_q[4] ),
    .X(_0018_));
 sky130_fd_sc_hd__clkbuf_4 _2589_ (.A(_0514_),
    .X(_0839_));
 sky130_fd_sc_hd__a32o_1 _2590_ (.A1(\usb2uart.u_usb_cdc.u_sie.phy_state_q[3] ),
    .A2(_2004_),
    .A3(_0591_),
    .B1(_0839_),
    .B2(\usb2uart.u_usb_cdc.u_sie.phy_state_q[9] ),
    .X(_0028_));
 sky130_fd_sc_hd__a21o_1 _2591_ (.A1(_2003_),
    .A2(_2004_),
    .B1(_0514_),
    .X(_0840_));
 sky130_fd_sc_hd__or2_2 _2592_ (.A(\usb2uart.u_usb_cdc.u_sie.phy_state_q[8] ),
    .B(\usb2uart.u_usb_cdc.u_sie.phy_state_q[2] ),
    .X(_0841_));
 sky130_fd_sc_hd__o211a_1 _2593_ (.A1(_0597_),
    .A2(_0836_),
    .B1(_0840_),
    .C1(_0841_),
    .X(_0027_));
 sky130_fd_sc_hd__nand2_1 _2594_ (.A(_2051_),
    .B(_2054_),
    .Y(_0842_));
 sky130_fd_sc_hd__nor2_1 _2595_ (.A(_0589_),
    .B(_0842_),
    .Y(_0843_));
 sky130_fd_sc_hd__buf_2 _2596_ (.A(\usb2uart.u_usb_cdc.u_sie.phy_state_q[7] ),
    .X(_0844_));
 sky130_fd_sc_hd__o21a_1 _2597_ (.A1(_0514_),
    .A2(_0843_),
    .B1(_0844_),
    .X(_0845_));
 sky130_fd_sc_hd__a31o_1 _2598_ (.A1(_2057_),
    .A2(_2056_),
    .A3(_0591_),
    .B1(_0845_),
    .X(_0026_));
 sky130_fd_sc_hd__a32o_1 _2599_ (.A1(\usb2uart.u_usb_cdc.u_sie.phy_state_q[0] ),
    .A2(_2004_),
    .A3(_0591_),
    .B1(_0514_),
    .B2(_0518_),
    .X(_0025_));
 sky130_fd_sc_hd__nand2_1 _2600_ (.A(_0521_),
    .B(\usb2uart.u_usb_cdc.u_sie.phy_state_q[6] ),
    .Y(_0846_));
 sky130_fd_sc_hd__o211a_1 _2601_ (.A1(_0552_),
    .A2(_0846_),
    .B1(_0595_),
    .C1(_0593_),
    .X(_0847_));
 sky130_fd_sc_hd__nor2_1 _2602_ (.A(_0514_),
    .B(_0847_),
    .Y(_0848_));
 sky130_fd_sc_hd__o21a_1 _2603_ (.A1(\usb2uart.u_usb_cdc.u_sie.phy_state_q[5] ),
    .A2(_0848_),
    .B1(_0840_),
    .X(_0024_));
 sky130_fd_sc_hd__nand2_1 _2604_ (.A(_2056_),
    .B(_0629_),
    .Y(_0849_));
 sky130_fd_sc_hd__a2bb2o_1 _2605_ (.A1_N(_2057_),
    .A2_N(_0849_),
    .B1(_0842_),
    .B2(_0844_),
    .X(_0850_));
 sky130_fd_sc_hd__a22o_1 _2606_ (.A1(\usb2uart.u_usb_cdc.u_sie.phy_state_q[4] ),
    .A2(_0515_),
    .B1(_0591_),
    .B2(_0850_),
    .X(_0023_));
 sky130_fd_sc_hd__and4bb_1 _2607_ (.A_N(_0719_),
    .B_N(\usb2uart.u_usb_cdc.u_ctrl_endp.class_q ),
    .C(_0718_),
    .D(_0762_),
    .X(_0851_));
 sky130_fd_sc_hd__nand2_1 _2608_ (.A(_2082_),
    .B(_0757_),
    .Y(_0852_));
 sky130_fd_sc_hd__and4b_1 _2609_ (.A_N(_0852_),
    .B(_2084_),
    .C(_2080_),
    .D(_0769_),
    .X(_0853_));
 sky130_fd_sc_hd__a31o_1 _2610_ (.A1(_0473_),
    .A2(_0681_),
    .A3(_0495_),
    .B1(_0853_),
    .X(_0854_));
 sky130_fd_sc_hd__o21a_1 _2611_ (.A1(_0695_),
    .A2(_0854_),
    .B1(\usb2uart.u_usb_cdc.u_ctrl_endp.req_q[5] ),
    .X(_0855_));
 sky130_fd_sc_hd__a21o_1 _2612_ (.A1(_0687_),
    .A2(_0851_),
    .B1(_0855_),
    .X(_0008_));
 sky130_fd_sc_hd__nand2_1 _2613_ (.A(_0492_),
    .B(_0457_),
    .Y(_0856_));
 sky130_fd_sc_hd__nor2_1 _2614_ (.A(_0856_),
    .B(_0707_),
    .Y(_0857_));
 sky130_fd_sc_hd__inv_2 _2615_ (.A(_0489_),
    .Y(_0858_));
 sky130_fd_sc_hd__and3_1 _2616_ (.A(_0687_),
    .B(_0688_),
    .C(_0858_),
    .X(_0859_));
 sky130_fd_sc_hd__o41a_1 _2617_ (.A1(_0859_),
    .A2(_0759_),
    .A3(_0698_),
    .A4(_0753_),
    .B1(\usb2uart.u_usb_cdc.u_ctrl_endp.req_q[0] ),
    .X(_0860_));
 sky130_fd_sc_hd__a31o_1 _2618_ (.A1(_2080_),
    .A2(_2082_),
    .A3(_0857_),
    .B1(_0860_),
    .X(_0001_));
 sky130_fd_sc_hd__nand2_1 _2619_ (.A(\usb2uart.u_usb_cdc.endp[0] ),
    .B(_2007_),
    .Y(_0861_));
 sky130_fd_sc_hd__or2_2 _2620_ (.A(_2077_),
    .B(_0861_),
    .X(_0862_));
 sky130_fd_sc_hd__inv_2 _2621_ (.A(_0862_),
    .Y(_0863_));
 sky130_fd_sc_hd__or2_1 _2622_ (.A(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_state_q[1] ),
    .B(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_full_o ),
    .X(_0864_));
 sky130_fd_sc_hd__and2b_1 _2623_ (.A_N(_0661_),
    .B(_0864_),
    .X(_0865_));
 sky130_fd_sc_hd__nor2_2 _2624_ (.A(_0862_),
    .B(_0865_),
    .Y(_0866_));
 sky130_fd_sc_hd__o21ba_1 _2625_ (.A1(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_state_q[1] ),
    .A2(_0863_),
    .B1_N(_0866_),
    .X(_0000_));
 sky130_fd_sc_hd__or3_1 _2626_ (.A(_0479_),
    .B(_0481_),
    .C(_0740_),
    .X(_0867_));
 sky130_fd_sc_hd__a22o_1 _2627_ (.A1(_0459_),
    .A2(_0711_),
    .B1(_0867_),
    .B2(\usb2uart.u_usb_cdc.u_ctrl_endp.req_q[4] ),
    .X(_0868_));
 sky130_fd_sc_hd__a22o_1 _2628_ (.A1(\usb2uart.u_usb_cdc.u_ctrl_endp.req_q[4] ),
    .A2(_0698_),
    .B1(_0868_),
    .B2(_2080_),
    .X(_0007_));
 sky130_fd_sc_hd__nor2_1 _2629_ (.A(_0714_),
    .B(_0730_),
    .Y(_0869_));
 sky130_fd_sc_hd__o31a_1 _2630_ (.A1(_0496_),
    .A2(_0695_),
    .A3(_0853_),
    .B1(\usb2uart.u_usb_cdc.u_ctrl_endp.req_q[3] ),
    .X(_0870_));
 sky130_fd_sc_hd__a21o_1 _2631_ (.A1(_0460_),
    .A2(_0869_),
    .B1(_0870_),
    .X(_0006_));
 sky130_fd_sc_hd__o21a_1 _2632_ (.A1(_0756_),
    .A2(_0758_),
    .B1(\usb2uart.u_usb_cdc.u_ctrl_endp.req_q[2] ),
    .X(_0871_));
 sky130_fd_sc_hd__a31o_1 _2633_ (.A1(\usb2uart.u_usb_cdc.u_ctrl_endp.req_q[9] ),
    .A2(_0759_),
    .A3(_0769_),
    .B1(_0871_),
    .X(_0005_));
 sky130_fd_sc_hd__o21a_1 _2634_ (.A1(_0792_),
    .A2(\usb2uart.u_usb_cdc.u_sie.u_phy_tx.data_q[0] ),
    .B1(\usb2uart.u_usb_cdc.u_sie.u_phy_tx.nrzi_q ),
    .X(\usb2uart.dp_tx ));
 sky130_fd_sc_hd__o21ba_1 _2635_ (.A1(_0792_),
    .A2(\usb2uart.u_usb_cdc.u_sie.u_phy_tx.data_q[0] ),
    .B1_N(\usb2uart.u_usb_cdc.u_sie.u_phy_tx.nrzi_q ),
    .X(\usb2uart.dn_tx ));
 sky130_fd_sc_hd__o41a_1 _2636_ (.A1(_0844_),
    .A2(_0553_),
    .A3(\usb2uart.u_usb_cdc.u_sie.phy_state_q[4] ),
    .A4(_0634_),
    .B1(_2003_),
    .X(_0872_));
 sky130_fd_sc_hd__o21ba_1 _2637_ (.A1(_0787_),
    .A2(_0872_),
    .B1_N(\usb2uart.u_usb_cdc.u_sie.u_phy_tx.clk_cnt_q[0] ),
    .X(_0042_));
 sky130_fd_sc_hd__or2_1 _2638_ (.A(\usb2uart.u_usb_cdc.u_sie.u_phy_tx.clk_cnt_q[1] ),
    .B(\usb2uart.u_usb_cdc.u_sie.u_phy_tx.clk_cnt_q[0] ),
    .X(_0873_));
 sky130_fd_sc_hd__o211a_1 _2639_ (.A1(_0787_),
    .A2(_0872_),
    .B1(_0873_),
    .C1(_0783_),
    .X(_0043_));
 sky130_fd_sc_hd__or2_1 _2640_ (.A(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.dn_q[0] ),
    .B(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.dn_q[1] ),
    .X(_0874_));
 sky130_fd_sc_hd__nand2_1 _2641_ (.A(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.dn_q[0] ),
    .B(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.dn_q[1] ),
    .Y(_0875_));
 sky130_fd_sc_hd__nand2_1 _2642_ (.A(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.dp_q[0] ),
    .B(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.dp_q[1] ),
    .Y(_0876_));
 sky130_fd_sc_hd__or2_1 _2643_ (.A(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.dp_q[0] ),
    .B(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.dp_q[1] ),
    .X(_0877_));
 sky130_fd_sc_hd__a22o_1 _2644_ (.A1(_0874_),
    .A2(_0875_),
    .B1(_0876_),
    .B2(_0877_),
    .X(_0878_));
 sky130_fd_sc_hd__nor2_1 _2645_ (.A(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.clk_cnt_q[0] ),
    .B(_0878_),
    .Y(_0040_));
 sky130_fd_sc_hd__or2b_1 _2646_ (.A(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.clk_cnt_q[0] ),
    .B_N(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.clk_cnt_q[1] ),
    .X(_0879_));
 sky130_fd_sc_hd__a21oi_1 _2647_ (.A1(_0795_),
    .A2(_0879_),
    .B1(_0878_),
    .Y(_0041_));
 sky130_fd_sc_hd__a21oi_1 _2648_ (.A1(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.rx_en_q ),
    .A2(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.cnt_q[5] ),
    .B1(\usb2uart.u_usb_cdc.u_ctrl_endp.usb_reset_q ),
    .Y(_0880_));
 sky130_fd_sc_hd__a21oi_1 _2649_ (.A1(\usb2uart.u_usb_cdc.u_ctrl_endp.usb_reset_q ),
    .A2(_0644_),
    .B1(_0880_),
    .Y(_0039_));
 sky130_fd_sc_hd__nor2_1 _2650_ (.A(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_state_q ),
    .B(_0779_),
    .Y(_0881_));
 sky130_fd_sc_hd__a31o_1 _2651_ (.A1(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_state_q ),
    .A2(_0487_),
    .A3(_0862_),
    .B1(_0881_),
    .X(_0038_));
 sky130_fd_sc_hd__or4_1 _2652_ (.A(\usb2uart.u_usb_cdc.endp[0] ),
    .B(\usb2uart.u_usb_cdc.endp[1] ),
    .C(\usb2uart.u_usb_cdc.endp[3] ),
    .D(\usb2uart.u_usb_cdc.endp[2] ),
    .X(_0882_));
 sky130_fd_sc_hd__buf_2 _2653_ (.A(_0882_),
    .X(_0883_));
 sky130_fd_sc_hd__or2_2 _2654_ (.A(_0589_),
    .B(_0777_),
    .X(_0884_));
 sky130_fd_sc_hd__nor2_1 _2655_ (.A(_0883_),
    .B(_0884_),
    .Y(\usb2uart.u_usb_cdc.ctrl_in_req ));
 sky130_fd_sc_hd__nand2_1 _2656_ (.A(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.rx_en_q ),
    .B(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.cnt_q[5] ),
    .Y(_0885_));
 sky130_fd_sc_hd__and2_1 _2657_ (.A(net58),
    .B(_0885_),
    .X(_0886_));
 sky130_fd_sc_hd__clkbuf_1 _2658_ (.A(_0886_),
    .X(\usb2uart.u_usb_cdc.u_bulk_endp.rstn ));
 sky130_fd_sc_hd__clkbuf_1 _2659_ (.A(net6),
    .X(_0887_));
 sky130_fd_sc_hd__clkbuf_1 _2660_ (.A(_0887_),
    .X(_2086_));
 sky130_fd_sc_hd__nand2_1 _2661_ (.A(_0521_),
    .B(_0527_),
    .Y(_0888_));
 sky130_fd_sc_hd__nor4_1 _2662_ (.A(_0517_),
    .B(_0519_),
    .C(_0551_),
    .D(_0888_),
    .Y(_0889_));
 sky130_fd_sc_hd__nand2_1 _2663_ (.A(\usb2uart.u_usb_cdc.u_sie.datain_toggle_q[0] ),
    .B(_2009_),
    .Y(_0890_));
 sky130_fd_sc_hd__o21a_1 _2664_ (.A1(\usb2uart.u_usb_cdc.u_sie.datain_toggle_q[0] ),
    .A2(_2009_),
    .B1(_0588_),
    .X(_0891_));
 sky130_fd_sc_hd__a31o_1 _2665_ (.A1(_0889_),
    .A2(_0890_),
    .A3(_0891_),
    .B1(\usb2uart.u_usb_cdc.u_sie.phy_state_q[9] ),
    .X(_0892_));
 sky130_fd_sc_hd__and3b_1 _2666_ (.A_N(_0533_),
    .B(_0531_),
    .C(\usb2uart.u_usb_cdc.u_sie.pid_q[2] ),
    .X(_0893_));
 sky130_fd_sc_hd__or4_1 _2667_ (.A(_2004_),
    .B(_0576_),
    .C(_0585_),
    .D(_0893_),
    .X(_0894_));
 sky130_fd_sc_hd__o21a_1 _2668_ (.A1(_0519_),
    .A2(_0551_),
    .B1(_2045_),
    .X(_0895_));
 sky130_fd_sc_hd__o31a_1 _2669_ (.A1(_0517_),
    .A2(_0888_),
    .A3(_0895_),
    .B1(_0518_),
    .X(_0896_));
 sky130_fd_sc_hd__and3_1 _2670_ (.A(\usb2uart.u_usb_cdc.u_sie.phy_state_q[9] ),
    .B(_0588_),
    .C(_0534_),
    .X(_0897_));
 sky130_fd_sc_hd__o32a_1 _2671_ (.A1(_0517_),
    .A2(_2045_),
    .A3(_0846_),
    .B1(_0518_),
    .B2(\usb2uart.u_usb_cdc.u_sie.phy_state_q[9] ),
    .X(_0898_));
 sky130_fd_sc_hd__or4b_1 _2672_ (.A(_0633_),
    .B(_0896_),
    .C(_0897_),
    .D_N(_0898_),
    .X(_0899_));
 sky130_fd_sc_hd__a21oi_1 _2673_ (.A1(\usb2uart.u_usb_cdc.u_sie.phy_state_q[9] ),
    .A2(_0894_),
    .B1(_0899_),
    .Y(_0900_));
 sky130_fd_sc_hd__mux2_1 _2674_ (.A0(\usb2uart.u_usb_cdc.u_sie.datain_toggle_q[0] ),
    .A1(_0892_),
    .S(_0900_),
    .X(_0901_));
 sky130_fd_sc_hd__clkbuf_1 _2675_ (.A(_0901_),
    .X(_0046_));
 sky130_fd_sc_hd__and3b_1 _2676_ (.A_N(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.cnt_q[5] ),
    .B(_0799_),
    .C(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.rx_en_q ),
    .X(_0902_));
 sky130_fd_sc_hd__a31o_1 _2677_ (.A1(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.rx_en_q ),
    .A2(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.cnt_q[5] ),
    .A3(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.cnt_q[2] ),
    .B1(_0902_),
    .X(_0903_));
 sky130_fd_sc_hd__nor2_2 _2678_ (.A(_2070_),
    .B(_0903_),
    .Y(_0904_));
 sky130_fd_sc_hd__buf_2 _2679_ (.A(_0904_),
    .X(_0905_));
 sky130_fd_sc_hd__inv_2 _2680_ (.A(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.cnt_q[2] ),
    .Y(_0906_));
 sky130_fd_sc_hd__o31ai_4 _2681_ (.A1(_0906_),
    .A2(_0799_),
    .A3(_0885_),
    .B1(_0825_),
    .Y(_0907_));
 sky130_fd_sc_hd__inv_2 _2682_ (.A(_0907_),
    .Y(_0908_));
 sky130_fd_sc_hd__and2_1 _2683_ (.A(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.cnt_q[0] ),
    .B(_0908_),
    .X(_0909_));
 sky130_fd_sc_hd__o21ba_1 _2684_ (.A1(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.cnt_q[0] ),
    .A2(_0905_),
    .B1_N(_0909_),
    .X(_0047_));
 sky130_fd_sc_hd__a21oi_1 _2685_ (.A1(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.cnt_q[0] ),
    .A2(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.cnt_q[1] ),
    .B1(_0903_),
    .Y(_0910_));
 sky130_fd_sc_hd__buf_2 _2686_ (.A(_0907_),
    .X(_0911_));
 sky130_fd_sc_hd__o22a_1 _2687_ (.A1(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.cnt_q[1] ),
    .A2(_0909_),
    .B1(_0910_),
    .B2(_0911_),
    .X(_0048_));
 sky130_fd_sc_hd__and3_1 _2688_ (.A(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.cnt_q[2] ),
    .B(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.cnt_q[0] ),
    .C(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.cnt_q[1] ),
    .X(_0912_));
 sky130_fd_sc_hd__and2_1 _2689_ (.A(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.cnt_q[3] ),
    .B(_0912_),
    .X(_0913_));
 sky130_fd_sc_hd__or2_1 _2690_ (.A(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.cnt_q[3] ),
    .B(_0912_),
    .X(_0914_));
 sky130_fd_sc_hd__and2b_1 _2691_ (.A_N(_0913_),
    .B(_0914_),
    .X(_0915_));
 sky130_fd_sc_hd__a22o_1 _2692_ (.A1(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.cnt_q[3] ),
    .A2(_0911_),
    .B1(_0905_),
    .B2(_0915_),
    .X(_0049_));
 sky130_fd_sc_hd__a21oi_1 _2693_ (.A1(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.cnt_q[4] ),
    .A2(_0913_),
    .B1(_0903_),
    .Y(_0916_));
 sky130_fd_sc_hd__a31o_1 _2694_ (.A1(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.cnt_q[3] ),
    .A2(_0908_),
    .A3(_0912_),
    .B1(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.cnt_q[4] ),
    .X(_0917_));
 sky130_fd_sc_hd__o21a_1 _2695_ (.A1(_0911_),
    .A2(_0916_),
    .B1(_0917_),
    .X(_0050_));
 sky130_fd_sc_hd__and3_1 _2696_ (.A(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.cnt_q[5] ),
    .B(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.cnt_q[4] ),
    .C(_0913_),
    .X(_0918_));
 sky130_fd_sc_hd__and2_1 _2697_ (.A(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.cnt_q[6] ),
    .B(_0918_),
    .X(_0919_));
 sky130_fd_sc_hd__o21ai_1 _2698_ (.A1(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.cnt_q[6] ),
    .A2(_0918_),
    .B1(_0905_),
    .Y(_0920_));
 sky130_fd_sc_hd__a2bb2o_1 _2699_ (.A1_N(_0919_),
    .A2_N(_0920_),
    .B1(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.cnt_q[6] ),
    .B2(_0911_),
    .X(_0051_));
 sky130_fd_sc_hd__and3_1 _2700_ (.A(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.cnt_q[6] ),
    .B(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.cnt_q[7] ),
    .C(_0918_),
    .X(_0921_));
 sky130_fd_sc_hd__o21ai_1 _2701_ (.A1(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.cnt_q[7] ),
    .A2(_0919_),
    .B1(_0904_),
    .Y(_0922_));
 sky130_fd_sc_hd__a2bb2o_1 _2702_ (.A1_N(_0921_),
    .A2_N(_0922_),
    .B1(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.cnt_q[7] ),
    .B2(_0911_),
    .X(_0052_));
 sky130_fd_sc_hd__nand2_1 _2703_ (.A(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.cnt_q[8] ),
    .B(_0921_),
    .Y(_0923_));
 sky130_fd_sc_hd__or2_1 _2704_ (.A(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.cnt_q[8] ),
    .B(_0921_),
    .X(_0924_));
 sky130_fd_sc_hd__a32o_1 _2705_ (.A1(_0905_),
    .A2(_0923_),
    .A3(_0924_),
    .B1(_0911_),
    .B2(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.cnt_q[8] ),
    .X(_0053_));
 sky130_fd_sc_hd__a21o_1 _2706_ (.A1(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.cnt_q[8] ),
    .A2(_0921_),
    .B1(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.cnt_q[9] ),
    .X(_0925_));
 sky130_fd_sc_hd__and3_1 _2707_ (.A(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.cnt_q[9] ),
    .B(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.cnt_q[8] ),
    .C(_0921_),
    .X(_0926_));
 sky130_fd_sc_hd__inv_2 _2708_ (.A(_0926_),
    .Y(_0927_));
 sky130_fd_sc_hd__a32o_1 _2709_ (.A1(_0905_),
    .A2(_0925_),
    .A3(_0927_),
    .B1(_0911_),
    .B2(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.cnt_q[9] ),
    .X(_0054_));
 sky130_fd_sc_hd__and2_1 _2710_ (.A(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.cnt_q[10] ),
    .B(_0926_),
    .X(_0928_));
 sky130_fd_sc_hd__o21ai_1 _2711_ (.A1(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.cnt_q[10] ),
    .A2(_0926_),
    .B1(_0904_),
    .Y(_0929_));
 sky130_fd_sc_hd__a2bb2o_1 _2712_ (.A1_N(_0928_),
    .A2_N(_0929_),
    .B1(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.cnt_q[10] ),
    .B2(_0911_),
    .X(_0055_));
 sky130_fd_sc_hd__nand2_1 _2713_ (.A(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.cnt_q[11] ),
    .B(_0928_),
    .Y(_0930_));
 sky130_fd_sc_hd__or2_1 _2714_ (.A(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.cnt_q[11] ),
    .B(_0928_),
    .X(_0931_));
 sky130_fd_sc_hd__a32o_1 _2715_ (.A1(_0905_),
    .A2(_0930_),
    .A3(_0931_),
    .B1(_0911_),
    .B2(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.cnt_q[11] ),
    .X(_0056_));
 sky130_fd_sc_hd__a31o_1 _2716_ (.A1(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.cnt_q[10] ),
    .A2(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.cnt_q[11] ),
    .A3(_0926_),
    .B1(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.cnt_q[12] ),
    .X(_0932_));
 sky130_fd_sc_hd__and3_1 _2717_ (.A(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.cnt_q[11] ),
    .B(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.cnt_q[12] ),
    .C(_0928_),
    .X(_0933_));
 sky130_fd_sc_hd__inv_2 _2718_ (.A(_0933_),
    .Y(_0934_));
 sky130_fd_sc_hd__a32o_1 _2719_ (.A1(_0905_),
    .A2(_0932_),
    .A3(_0934_),
    .B1(_0911_),
    .B2(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.cnt_q[12] ),
    .X(_0057_));
 sky130_fd_sc_hd__or2_1 _2720_ (.A(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.cnt_q[13] ),
    .B(_0933_),
    .X(_0935_));
 sky130_fd_sc_hd__and2_1 _2721_ (.A(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.cnt_q[13] ),
    .B(_0933_),
    .X(_0936_));
 sky130_fd_sc_hd__inv_2 _2722_ (.A(_0936_),
    .Y(_0937_));
 sky130_fd_sc_hd__a32o_1 _2723_ (.A1(_0905_),
    .A2(_0935_),
    .A3(_0937_),
    .B1(_0907_),
    .B2(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.cnt_q[13] ),
    .X(_0058_));
 sky130_fd_sc_hd__nand2_1 _2724_ (.A(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.cnt_q[14] ),
    .B(_0936_),
    .Y(_0938_));
 sky130_fd_sc_hd__or2_1 _2725_ (.A(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.cnt_q[14] ),
    .B(_0936_),
    .X(_0939_));
 sky130_fd_sc_hd__a32o_1 _2726_ (.A1(_0905_),
    .A2(_0938_),
    .A3(_0939_),
    .B1(_0907_),
    .B2(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.cnt_q[14] ),
    .X(_0059_));
 sky130_fd_sc_hd__a31o_1 _2727_ (.A1(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.cnt_q[13] ),
    .A2(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.cnt_q[14] ),
    .A3(_0933_),
    .B1(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.cnt_q[15] ),
    .X(_0940_));
 sky130_fd_sc_hd__and3_1 _2728_ (.A(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.cnt_q[14] ),
    .B(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.cnt_q[15] ),
    .C(_0936_),
    .X(_0941_));
 sky130_fd_sc_hd__inv_2 _2729_ (.A(_0941_),
    .Y(_0942_));
 sky130_fd_sc_hd__a32o_1 _2730_ (.A1(_0905_),
    .A2(_0940_),
    .A3(_0942_),
    .B1(_0907_),
    .B2(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.cnt_q[15] ),
    .X(_0060_));
 sky130_fd_sc_hd__a21o_1 _2731_ (.A1(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.cnt_q[16] ),
    .A2(_0941_),
    .B1(_0903_),
    .X(_0943_));
 sky130_fd_sc_hd__nand2_1 _2732_ (.A(_0908_),
    .B(_0943_),
    .Y(_0944_));
 sky130_fd_sc_hd__a21o_1 _2733_ (.A1(_0904_),
    .A2(_0941_),
    .B1(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.cnt_q[16] ),
    .X(_0945_));
 sky130_fd_sc_hd__and2_1 _2734_ (.A(_0944_),
    .B(_0945_),
    .X(_0946_));
 sky130_fd_sc_hd__clkbuf_1 _2735_ (.A(_0946_),
    .X(_0061_));
 sky130_fd_sc_hd__and3_1 _2736_ (.A(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.cnt_q[16] ),
    .B(_0904_),
    .C(_0941_),
    .X(_0947_));
 sky130_fd_sc_hd__mux2_1 _2737_ (.A0(_0947_),
    .A1(_0944_),
    .S(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.cnt_q[17] ),
    .X(_0948_));
 sky130_fd_sc_hd__clkbuf_1 _2738_ (.A(_0948_),
    .X(_0062_));
 sky130_fd_sc_hd__mux2_1 _2739_ (.A0(_0872_),
    .A1(_0781_),
    .S(_0783_),
    .X(_0949_));
 sky130_fd_sc_hd__clkbuf_1 _2740_ (.A(_0949_),
    .X(_0063_));
 sky130_fd_sc_hd__inv_2 _2741_ (.A(net4),
    .Y(_0950_));
 sky130_fd_sc_hd__clkbuf_4 _2742_ (.A(_0950_),
    .X(_0044_));
 sky130_fd_sc_hd__clkbuf_4 _2743_ (.A(net4),
    .X(_0951_));
 sky130_fd_sc_hd__inv_2 _2744_ (.A(_0951_),
    .Y(_0045_));
 sky130_fd_sc_hd__a21o_1 _2745_ (.A1(\usb2uart.u_usb_cdc.u_sie.u_phy_tx.tx_state_q[2] ),
    .A2(_0790_),
    .B1(\usb2uart.u_usb_cdc.u_sie.u_phy_tx.tx_state_q[1] ),
    .X(_0952_));
 sky130_fd_sc_hd__a31o_1 _2746_ (.A1(\usb2uart.u_usb_cdc.u_sie.u_phy_tx.tx_state_q[3] ),
    .A2(\usb2uart.u_usb_cdc.u_sie.u_phy_tx.data_q[1] ),
    .A3(_0785_),
    .B1(_0952_),
    .X(_0953_));
 sky130_fd_sc_hd__nor2_1 _2747_ (.A(_0589_),
    .B(_2063_),
    .Y(_0954_));
 sky130_fd_sc_hd__inv_2 _2748_ (.A(\usb2uart.u_usb_cdc.u_sie.crc16_q[7] ),
    .Y(_0955_));
 sky130_fd_sc_hd__a22o_1 _2749_ (.A1(\usb2uart.u_usb_cdc.u_sie.pid_q[0] ),
    .A2(\usb2uart.u_usb_cdc.u_sie.phy_state_q[11] ),
    .B1(\usb2uart.u_usb_cdc.u_sie.phy_state_q[10] ),
    .B2(_0955_),
    .X(_0956_));
 sky130_fd_sc_hd__inv_2 _2750_ (.A(\usb2uart.u_usb_cdc.u_sie.phy_state_q[4] ),
    .Y(_0957_));
 sky130_fd_sc_hd__a2bb2o_1 _2751_ (.A1_N(\usb2uart.u_usb_cdc.u_sie.crc16_q[15] ),
    .A2_N(_0957_),
    .B1(\usb2uart.u_usb_cdc.u_sie.phy_state_q[7] ),
    .B2(_0517_),
    .X(_0958_));
 sky130_fd_sc_hd__or3b_1 _2752_ (.A(_0956_),
    .B(_0958_),
    .C_N(_0849_),
    .X(_0959_));
 sky130_fd_sc_hd__a221o_1 _2753_ (.A1(\usb2uart.u_usb_cdc.u_sie.u_phy_tx.data_q[1] ),
    .A2(_0785_),
    .B1(_0954_),
    .B2(_0959_),
    .C1(_0782_),
    .X(_0960_));
 sky130_fd_sc_hd__nor2_1 _2754_ (.A(\usb2uart.u_usb_cdc.u_sie.u_phy_tx.tx_state_q[1] ),
    .B(_0794_),
    .Y(_0961_));
 sky130_fd_sc_hd__a21o_1 _2755_ (.A1(_0953_),
    .A2(_0960_),
    .B1(_0961_),
    .X(_0962_));
 sky130_fd_sc_hd__or2_1 _2756_ (.A(\usb2uart.u_usb_cdc.u_sie.u_phy_tx.tx_state_q[1] ),
    .B(_0794_),
    .X(_0963_));
 sky130_fd_sc_hd__or2_1 _2757_ (.A(\usb2uart.u_usb_cdc.u_sie.u_phy_tx.data_q[1] ),
    .B(_0963_),
    .X(_0964_));
 sky130_fd_sc_hd__or2_1 _2758_ (.A(_0781_),
    .B(_0963_),
    .X(_0965_));
 sky130_fd_sc_hd__and2_1 _2759_ (.A(_0780_),
    .B(_0965_),
    .X(_0966_));
 sky130_fd_sc_hd__a32o_1 _2760_ (.A1(_0962_),
    .A2(_0964_),
    .A3(_0966_),
    .B1(_0788_),
    .B2(\usb2uart.u_usb_cdc.u_sie.u_phy_tx.data_q[0] ),
    .X(_0064_));
 sky130_fd_sc_hd__o21a_1 _2761_ (.A1(_0785_),
    .A2(_0961_),
    .B1(_0965_),
    .X(_0967_));
 sky130_fd_sc_hd__and3_1 _2762_ (.A(_0781_),
    .B(_0791_),
    .C(_0954_),
    .X(_0968_));
 sky130_fd_sc_hd__inv_2 _2763_ (.A(\usb2uart.u_usb_cdc.u_sie.crc16_q[6] ),
    .Y(_0969_));
 sky130_fd_sc_hd__nor2_1 _2764_ (.A(\usb2uart.u_usb_cdc.u_sie.crc16_q[14] ),
    .B(_0957_),
    .Y(_0970_));
 sky130_fd_sc_hd__a221o_1 _2765_ (.A1(_0844_),
    .A2(_0521_),
    .B1(\usb2uart.u_usb_cdc.u_sie.phy_state_q[11] ),
    .B2(\usb2uart.u_usb_cdc.u_sie.pid_q[1] ),
    .C1(_0970_),
    .X(_0971_));
 sky130_fd_sc_hd__a211o_1 _2766_ (.A1(\usb2uart.u_usb_cdc.u_sie.phy_state_q[10] ),
    .A2(_0969_),
    .B1(_0971_),
    .C1(_0553_),
    .X(_0972_));
 sky130_fd_sc_hd__a221o_1 _2767_ (.A1(\usb2uart.u_usb_cdc.u_sie.u_phy_tx.data_q[2] ),
    .A2(_0967_),
    .B1(_0968_),
    .B2(_0972_),
    .C1(_0788_),
    .X(_0973_));
 sky130_fd_sc_hd__o21a_1 _2768_ (.A1(\usb2uart.u_usb_cdc.u_sie.u_phy_tx.data_q[1] ),
    .A2(_0780_),
    .B1(_0973_),
    .X(_0065_));
 sky130_fd_sc_hd__inv_2 _2769_ (.A(\usb2uart.u_usb_cdc.u_sie.phy_state_q[10] ),
    .Y(_0974_));
 sky130_fd_sc_hd__o2bb2a_1 _2770_ (.A1_N(_0844_),
    .A2_N(\usb2uart.u_usb_cdc.u_sie.data_q[2] ),
    .B1(_0974_),
    .B2(\usb2uart.u_usb_cdc.u_sie.crc16_q[5] ),
    .X(_0975_));
 sky130_fd_sc_hd__o22a_1 _2771_ (.A1(_0532_),
    .A2(_0835_),
    .B1(\usb2uart.u_usb_cdc.u_sie.crc16_q[13] ),
    .B2(_0957_),
    .X(_0976_));
 sky130_fd_sc_hd__o211ai_1 _2772_ (.A1(_0630_),
    .A2(_2055_),
    .B1(_0975_),
    .C1(_0976_),
    .Y(_0977_));
 sky130_fd_sc_hd__a221o_1 _2773_ (.A1(\usb2uart.u_usb_cdc.u_sie.u_phy_tx.data_q[3] ),
    .A2(_0967_),
    .B1(_0968_),
    .B2(_0977_),
    .C1(_0784_),
    .X(_0978_));
 sky130_fd_sc_hd__o21a_1 _2774_ (.A1(\usb2uart.u_usb_cdc.u_sie.u_phy_tx.data_q[2] ),
    .A2(_0780_),
    .B1(_0978_),
    .X(_0066_));
 sky130_fd_sc_hd__mux2_2 _2775_ (.A0(\usb2uart.u_usb_cdc.u_sie.datain_toggle_q[0] ),
    .A1(\usb2uart.u_usb_cdc.u_sie.datain_toggle_q[1] ),
    .S(\usb2uart.u_usb_cdc.endp[0] ),
    .X(_0979_));
 sky130_fd_sc_hd__inv_2 _2776_ (.A(\usb2uart.u_usb_cdc.u_sie.crc16_q[12] ),
    .Y(_0980_));
 sky130_fd_sc_hd__a2bb2o_1 _2777_ (.A1_N(_0974_),
    .A2_N(\usb2uart.u_usb_cdc.u_sie.crc16_q[4] ),
    .B1(\usb2uart.u_usb_cdc.u_sie.phy_state_q[7] ),
    .B2(_0519_),
    .X(_0981_));
 sky130_fd_sc_hd__a221o_1 _2778_ (.A1(\usb2uart.u_usb_cdc.u_sie.pid_q[3] ),
    .A2(\usb2uart.u_usb_cdc.u_sie.phy_state_q[11] ),
    .B1(_0980_),
    .B2(\usb2uart.u_usb_cdc.u_sie.phy_state_q[4] ),
    .C1(_0981_),
    .X(_0982_));
 sky130_fd_sc_hd__a211o_1 _2779_ (.A1(_0553_),
    .A2(_0979_),
    .B1(_0982_),
    .C1(_0631_),
    .X(_0983_));
 sky130_fd_sc_hd__a221o_1 _2780_ (.A1(\usb2uart.u_usb_cdc.u_sie.u_phy_tx.data_q[4] ),
    .A2(_2063_),
    .B1(_0954_),
    .B2(_0983_),
    .C1(_0782_),
    .X(_0984_));
 sky130_fd_sc_hd__a32o_1 _2781_ (.A1(\usb2uart.u_usb_cdc.u_sie.u_phy_tx.tx_state_q[3] ),
    .A2(\usb2uart.u_usb_cdc.u_sie.u_phy_tx.data_q[4] ),
    .A3(_0785_),
    .B1(_0952_),
    .B2(_0984_),
    .X(_0985_));
 sky130_fd_sc_hd__or2_1 _2782_ (.A(_0961_),
    .B(_0985_),
    .X(_0986_));
 sky130_fd_sc_hd__or2_1 _2783_ (.A(\usb2uart.u_usb_cdc.u_sie.u_phy_tx.data_q[4] ),
    .B(_0963_),
    .X(_0987_));
 sky130_fd_sc_hd__a32o_1 _2784_ (.A1(_0966_),
    .A2(_0986_),
    .A3(_0987_),
    .B1(_0788_),
    .B2(\usb2uart.u_usb_cdc.u_sie.u_phy_tx.data_q[3] ),
    .X(_0067_));
 sky130_fd_sc_hd__a2bb2o_1 _2785_ (.A1_N(\usb2uart.u_usb_cdc.u_sie.crc16_q[11] ),
    .A2_N(_0957_),
    .B1(\usb2uart.u_usb_cdc.u_sie.phy_state_q[7] ),
    .B2(\usb2uart.u_usb_cdc.u_sie.data_q[4] ),
    .X(_0988_));
 sky130_fd_sc_hd__o22a_1 _2786_ (.A1(\usb2uart.u_usb_cdc.u_sie.pid_q[0] ),
    .A2(_0835_),
    .B1(_0974_),
    .B2(\usb2uart.u_usb_cdc.u_sie.crc16_q[3] ),
    .X(_0989_));
 sky130_fd_sc_hd__or3b_1 _2787_ (.A(_0988_),
    .B(_0631_),
    .C_N(_0989_),
    .X(_0990_));
 sky130_fd_sc_hd__a221o_1 _2788_ (.A1(\usb2uart.u_usb_cdc.u_sie.u_phy_tx.data_q[5] ),
    .A2(_0785_),
    .B1(_0954_),
    .B2(_0990_),
    .C1(_0782_),
    .X(_0991_));
 sky130_fd_sc_hd__a31o_1 _2789_ (.A1(\usb2uart.u_usb_cdc.u_sie.u_phy_tx.tx_state_q[3] ),
    .A2(\usb2uart.u_usb_cdc.u_sie.u_phy_tx.data_q[5] ),
    .A3(_0785_),
    .B1(_0961_),
    .X(_0992_));
 sky130_fd_sc_hd__a21o_1 _2790_ (.A1(_0952_),
    .A2(_0991_),
    .B1(_0992_),
    .X(_0993_));
 sky130_fd_sc_hd__or2_1 _2791_ (.A(\usb2uart.u_usb_cdc.u_sie.u_phy_tx.data_q[5] ),
    .B(_0963_),
    .X(_0994_));
 sky130_fd_sc_hd__a32o_1 _2792_ (.A1(_0966_),
    .A2(_0993_),
    .A3(_0994_),
    .B1(_0788_),
    .B2(\usb2uart.u_usb_cdc.u_sie.u_phy_tx.data_q[4] ),
    .X(_0068_));
 sky130_fd_sc_hd__o2bb2a_1 _2793_ (.A1_N(\usb2uart.u_usb_cdc.u_sie.phy_state_q[7] ),
    .A2_N(\usb2uart.u_usb_cdc.u_sie.data_q[5] ),
    .B1(_0974_),
    .B2(\usb2uart.u_usb_cdc.u_sie.crc16_q[2] ),
    .X(_0995_));
 sky130_fd_sc_hd__o221a_1 _2794_ (.A1(\usb2uart.u_usb_cdc.u_sie.pid_q[1] ),
    .A2(_0835_),
    .B1(\usb2uart.u_usb_cdc.u_sie.crc16_q[10] ),
    .B2(_0957_),
    .C1(_0995_),
    .X(_0996_));
 sky130_fd_sc_hd__o21ai_1 _2795_ (.A1(_0589_),
    .A2(_0996_),
    .B1(_0781_),
    .Y(_0997_));
 sky130_fd_sc_hd__a21oi_1 _2796_ (.A1(_0781_),
    .A2(\usb2uart.u_usb_cdc.u_sie.u_phy_tx.tx_state_q[2] ),
    .B1(\usb2uart.u_usb_cdc.u_sie.u_phy_tx.tx_state_q[1] ),
    .Y(_0998_));
 sky130_fd_sc_hd__nor2_1 _2797_ (.A(_0785_),
    .B(_0998_),
    .Y(_0999_));
 sky130_fd_sc_hd__a221o_1 _2798_ (.A1(\usb2uart.u_usb_cdc.u_sie.u_phy_tx.data_q[6] ),
    .A2(_0967_),
    .B1(_0997_),
    .B2(_0999_),
    .C1(_0784_),
    .X(_1000_));
 sky130_fd_sc_hd__o21a_1 _2799_ (.A1(\usb2uart.u_usb_cdc.u_sie.u_phy_tx.data_q[5] ),
    .A2(_0780_),
    .B1(_1000_),
    .X(_0069_));
 sky130_fd_sc_hd__inv_2 _2800_ (.A(\usb2uart.u_usb_cdc.u_sie.crc16_q[9] ),
    .Y(_1001_));
 sky130_fd_sc_hd__a221o_1 _2801_ (.A1(_0532_),
    .A2(\usb2uart.u_usb_cdc.u_sie.phy_state_q[11] ),
    .B1(_1001_),
    .B2(\usb2uart.u_usb_cdc.u_sie.phy_state_q[4] ),
    .C1(_2056_),
    .X(_1002_));
 sky130_fd_sc_hd__a221o_1 _2802_ (.A1(_0844_),
    .A2(\usb2uart.u_usb_cdc.u_sie.data_q[6] ),
    .B1(\usb2uart.u_usb_cdc.u_sie.phy_state_q[10] ),
    .B2(_0619_),
    .C1(_1002_),
    .X(_1003_));
 sky130_fd_sc_hd__a21bo_1 _2803_ (.A1(_2003_),
    .A2(_1003_),
    .B1_N(_0781_),
    .X(_1004_));
 sky130_fd_sc_hd__a221o_1 _2804_ (.A1(\usb2uart.u_usb_cdc.u_sie.u_phy_tx.data_q[7] ),
    .A2(_0967_),
    .B1(_0999_),
    .B2(_1004_),
    .C1(_0784_),
    .X(_1005_));
 sky130_fd_sc_hd__o21a_1 _2805_ (.A1(\usb2uart.u_usb_cdc.u_sie.u_phy_tx.data_q[6] ),
    .A2(_0780_),
    .B1(_1005_),
    .X(_0070_));
 sky130_fd_sc_hd__o2bb2a_1 _2806_ (.A1_N(_0844_),
    .A2_N(\usb2uart.u_usb_cdc.u_sie.data_q[7] ),
    .B1(_0835_),
    .B2(\usb2uart.u_usb_cdc.u_sie.pid_q[3] ),
    .X(_1006_));
 sky130_fd_sc_hd__o221a_1 _2807_ (.A1(_0974_),
    .A2(\usb2uart.u_usb_cdc.u_sie.crc16_q[0] ),
    .B1(_0957_),
    .B2(\usb2uart.u_usb_cdc.u_sie.crc16_q[8] ),
    .C1(_1006_),
    .X(_1007_));
 sky130_fd_sc_hd__o21ai_1 _2808_ (.A1(_0849_),
    .A2(_0979_),
    .B1(_1007_),
    .Y(_1008_));
 sky130_fd_sc_hd__a31o_1 _2809_ (.A1(_0791_),
    .A2(_0872_),
    .A3(_1008_),
    .B1(_0793_),
    .X(_1009_));
 sky130_fd_sc_hd__nor2_1 _2810_ (.A(_0788_),
    .B(_0967_),
    .Y(_1010_));
 sky130_fd_sc_hd__a22o_1 _2811_ (.A1(\usb2uart.u_usb_cdc.u_sie.u_phy_tx.data_q[7] ),
    .A2(_0788_),
    .B1(_1009_),
    .B2(_1010_),
    .X(_0071_));
 sky130_fd_sc_hd__a21oi_1 _2812_ (.A1(\usb2uart.u_usb_cdc.u_sie.u_phy_tx.bit_cnt_q[0] ),
    .A2(_0965_),
    .B1(_0788_),
    .Y(_1011_));
 sky130_fd_sc_hd__a21o_1 _2813_ (.A1(\usb2uart.u_usb_cdc.u_sie.u_phy_tx.bit_cnt_q[0] ),
    .A2(_0788_),
    .B1(_1011_),
    .X(_0072_));
 sky130_fd_sc_hd__nand2_1 _2814_ (.A(_0780_),
    .B(_0965_),
    .Y(_1012_));
 sky130_fd_sc_hd__or3b_1 _2815_ (.A(_1012_),
    .B(\usb2uart.u_usb_cdc.u_sie.u_phy_tx.bit_cnt_q[0] ),
    .C_N(\usb2uart.u_usb_cdc.u_sie.u_phy_tx.bit_cnt_q[1] ),
    .X(_1013_));
 sky130_fd_sc_hd__o21a_1 _2816_ (.A1(\usb2uart.u_usb_cdc.u_sie.u_phy_tx.bit_cnt_q[1] ),
    .A2(_1011_),
    .B1(_1013_),
    .X(_0073_));
 sky130_fd_sc_hd__o21a_1 _2817_ (.A1(\usb2uart.u_usb_cdc.u_sie.u_phy_tx.bit_cnt_q[0] ),
    .A2(\usb2uart.u_usb_cdc.u_sie.u_phy_tx.bit_cnt_q[1] ),
    .B1(\usb2uart.u_usb_cdc.u_sie.u_phy_tx.bit_cnt_q[2] ),
    .X(_1014_));
 sky130_fd_sc_hd__o21ba_1 _2818_ (.A1(_0781_),
    .A2(_0794_),
    .B1_N(_0785_),
    .X(_1015_));
 sky130_fd_sc_hd__o32a_1 _2819_ (.A1(_1012_),
    .A2(_1014_),
    .A3(_1015_),
    .B1(_0780_),
    .B2(\usb2uart.u_usb_cdc.u_sie.u_phy_tx.bit_cnt_q[2] ),
    .X(_0074_));
 sky130_fd_sc_hd__a21o_1 _2820_ (.A1(\usb2uart.u_usb_cdc.u_sie.u_phy_tx.data_q[0] ),
    .A2(_2060_),
    .B1(_0783_),
    .X(_1016_));
 sky130_fd_sc_hd__nor2_1 _2821_ (.A(_0781_),
    .B(_0791_),
    .Y(_1017_));
 sky130_fd_sc_hd__a211o_1 _2822_ (.A1(\usb2uart.u_usb_cdc.u_sie.u_phy_tx.tx_state_q[2] ),
    .A2(_0782_),
    .B1(_1017_),
    .C1(\usb2uart.u_usb_cdc.u_sie.u_phy_tx.tx_state_q[3] ),
    .X(_1018_));
 sky130_fd_sc_hd__a22o_1 _2823_ (.A1(_0780_),
    .A2(_1018_),
    .B1(_1016_),
    .B2(\usb2uart.u_usb_cdc.u_sie.u_phy_tx.nrzi_q ),
    .X(_1019_));
 sky130_fd_sc_hd__o21bai_1 _2824_ (.A1(\usb2uart.u_usb_cdc.u_sie.u_phy_tx.nrzi_q ),
    .A2(_1016_),
    .B1_N(_1019_),
    .Y(_0075_));
 sky130_fd_sc_hd__a31o_1 _2825_ (.A1(_0787_),
    .A2(_0792_),
    .A3(_0790_),
    .B1(\usb2uart.u_usb_cdc.u_sie.u_phy_tx.tx_state_q[1] ),
    .X(_1020_));
 sky130_fd_sc_hd__and3_1 _2826_ (.A(\usb2uart.u_usb_cdc.u_sie.u_phy_tx.data_q[0] ),
    .B(_0780_),
    .C(_1020_),
    .X(_1021_));
 sky130_fd_sc_hd__mux2_1 _2827_ (.A0(_1021_),
    .A1(_0783_),
    .S(\usb2uart.u_usb_cdc.u_sie.u_phy_tx.stuffing_cnt_q[0] ),
    .X(_1022_));
 sky130_fd_sc_hd__clkbuf_1 _2828_ (.A(_1022_),
    .X(_0076_));
 sky130_fd_sc_hd__or2_1 _2829_ (.A(\usb2uart.u_usb_cdc.u_sie.u_phy_tx.stuffing_cnt_q[0] ),
    .B(\usb2uart.u_usb_cdc.u_sie.u_phy_tx.stuffing_cnt_q[1] ),
    .X(_1023_));
 sky130_fd_sc_hd__nand2_1 _2830_ (.A(\usb2uart.u_usb_cdc.u_sie.u_phy_tx.stuffing_cnt_q[0] ),
    .B(\usb2uart.u_usb_cdc.u_sie.u_phy_tx.stuffing_cnt_q[1] ),
    .Y(_1024_));
 sky130_fd_sc_hd__a32o_1 _2831_ (.A1(_1021_),
    .A2(_1023_),
    .A3(_1024_),
    .B1(_0783_),
    .B2(\usb2uart.u_usb_cdc.u_sie.u_phy_tx.stuffing_cnt_q[1] ),
    .X(_0077_));
 sky130_fd_sc_hd__a41o_1 _2832_ (.A1(\usb2uart.u_usb_cdc.u_sie.u_phy_tx.clk_cnt_q[1] ),
    .A2(\usb2uart.u_usb_cdc.u_sie.u_phy_tx.clk_cnt_q[0] ),
    .A3(\usb2uart.u_usb_cdc.u_sie.u_phy_tx.stuffing_cnt_q[0] ),
    .A4(\usb2uart.u_usb_cdc.u_sie.u_phy_tx.stuffing_cnt_q[1] ),
    .B1(\usb2uart.u_usb_cdc.u_sie.u_phy_tx.stuffing_cnt_q[2] ),
    .X(_1025_));
 sky130_fd_sc_hd__a31o_1 _2833_ (.A1(\usb2uart.u_usb_cdc.u_sie.u_phy_tx.data_q[0] ),
    .A2(_2059_),
    .A3(_1020_),
    .B1(_0783_),
    .X(_1026_));
 sky130_fd_sc_hd__and2_1 _2834_ (.A(_1025_),
    .B(_1026_),
    .X(_1027_));
 sky130_fd_sc_hd__clkbuf_1 _2835_ (.A(_1027_),
    .X(_0078_));
 sky130_fd_sc_hd__and3_1 _2836_ (.A(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.cnt_q[16] ),
    .B(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.cnt_q[17] ),
    .C(_0826_),
    .X(_1028_));
 sky130_fd_sc_hd__a31o_1 _2837_ (.A1(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.cnt_q[9] ),
    .A2(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.cnt_q[8] ),
    .A3(_1028_),
    .B1(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.rx_en_q ),
    .X(_0079_));
 sky130_fd_sc_hd__a32o_1 _2838_ (.A1(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.cnt_q[0] ),
    .A2(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.cnt_q[1] ),
    .A3(_0885_),
    .B1(_0799_),
    .B2(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.rx_en_q ),
    .X(_1029_));
 sky130_fd_sc_hd__a21oi_1 _2839_ (.A1(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.cnt_q[2] ),
    .A2(_1029_),
    .B1(_0902_),
    .Y(_1030_));
 sky130_fd_sc_hd__a31o_1 _2840_ (.A1(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.cnt_q[0] ),
    .A2(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.cnt_q[1] ),
    .A3(_0826_),
    .B1(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.cnt_q[2] ),
    .X(_1031_));
 sky130_fd_sc_hd__o21a_1 _2841_ (.A1(_0795_),
    .A2(_1030_),
    .B1(_1031_),
    .X(_0080_));
 sky130_fd_sc_hd__and2b_1 _2842_ (.A_N(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.rx_en_q ),
    .B(_0918_),
    .X(_1032_));
 sky130_fd_sc_hd__a31o_1 _2843_ (.A1(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.rx_en_q ),
    .A2(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.cnt_q[2] ),
    .A3(_0799_),
    .B1(_1032_),
    .X(_1033_));
 sky130_fd_sc_hd__and3_1 _2844_ (.A(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.cnt_q[4] ),
    .B(_0826_),
    .C(_0913_),
    .X(_1034_));
 sky130_fd_sc_hd__o2bb2a_1 _2845_ (.A1_N(_0826_),
    .A2_N(_1033_),
    .B1(_1034_),
    .B2(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.cnt_q[5] ),
    .X(_0081_));
 sky130_fd_sc_hd__o21ai_1 _2846_ (.A1(_0819_),
    .A2(_0821_),
    .B1(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.rx_state_q[2] ),
    .Y(_1035_));
 sky130_fd_sc_hd__o31ai_1 _2847_ (.A1(_0819_),
    .A2(_0820_),
    .A3(_1035_),
    .B1(_0826_),
    .Y(_1036_));
 sky130_fd_sc_hd__and2_1 _2848_ (.A(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.rx_state_q[2] ),
    .B(_0823_),
    .X(_1037_));
 sky130_fd_sc_hd__or3_1 _2849_ (.A(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.rx_state_q[0] ),
    .B(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.rx_state_q[3] ),
    .C(_2068_),
    .X(_1038_));
 sky130_fd_sc_hd__o32a_1 _2850_ (.A1(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.dn_q[0] ),
    .A2(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.dp_q[0] ),
    .A3(_2066_),
    .B1(_1037_),
    .B2(_1038_),
    .X(_1039_));
 sky130_fd_sc_hd__a211o_1 _2851_ (.A1(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.rx_state_q[2] ),
    .A2(_0801_),
    .B1(_1036_),
    .C1(_1039_),
    .X(_1040_));
 sky130_fd_sc_hd__mux2_1 _2852_ (.A0(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.rx_valid_fd ),
    .A1(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.rx_valid_fq ),
    .S(_1040_),
    .X(_1041_));
 sky130_fd_sc_hd__clkbuf_1 _2853_ (.A(_1041_),
    .X(_0082_));
 sky130_fd_sc_hd__or3_1 _2854_ (.A(_2070_),
    .B(_0810_),
    .C(_0817_),
    .X(_1042_));
 sky130_fd_sc_hd__xnor2_1 _2855_ (.A(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.rx_valid_fd ),
    .B(_1042_),
    .Y(_0083_));
 sky130_fd_sc_hd__or2_1 _2856_ (.A(net7),
    .B(_1028_),
    .X(_1043_));
 sky130_fd_sc_hd__clkbuf_1 _2857_ (.A(_1043_),
    .X(_0084_));
 sky130_fd_sc_hd__nor4_1 _2858_ (.A(_0593_),
    .B(_0534_),
    .C(_0576_),
    .D(_0585_),
    .Y(_1044_));
 sky130_fd_sc_hd__a21oi_1 _2859_ (.A1(_0597_),
    .A2(_0593_),
    .B1(_1044_),
    .Y(_1045_));
 sky130_fd_sc_hd__or4_1 _2860_ (.A(_2004_),
    .B(_0633_),
    .C(_0627_),
    .D(_1045_),
    .X(_1046_));
 sky130_fd_sc_hd__inv_2 _2861_ (.A(\usb2uart.u_usb_cdc.u_sie.dataout_toggle_q[0] ),
    .Y(_1047_));
 sky130_fd_sc_hd__mux2_1 _2862_ (.A0(\usb2uart.u_usb_cdc.u_sie.dataout_toggle_q[0] ),
    .A1(\usb2uart.u_usb_cdc.u_sie.dataout_toggle_q[1] ),
    .S(\usb2uart.u_usb_cdc.endp[0] ),
    .X(_1048_));
 sky130_fd_sc_hd__xnor2_1 _2863_ (.A(\usb2uart.u_usb_cdc.u_sie.pid_q[3] ),
    .B(_1048_),
    .Y(_1049_));
 sky130_fd_sc_hd__nand2_1 _2864_ (.A(_2007_),
    .B(_1049_),
    .Y(_1050_));
 sky130_fd_sc_hd__nand2_1 _2865_ (.A(_0623_),
    .B(_0622_),
    .Y(_1051_));
 sky130_fd_sc_hd__or4_1 _2866_ (.A(_0606_),
    .B(_0620_),
    .C(_0617_),
    .D(_1051_),
    .X(_1052_));
 sky130_fd_sc_hd__or4_1 _2867_ (.A(_0601_),
    .B(_0614_),
    .C(_0621_),
    .D(_1052_),
    .X(_1053_));
 sky130_fd_sc_hd__or4_2 _2868_ (.A(\usb2uart.u_usb_cdc.u_sie.crc16_q[7] ),
    .B(_0613_),
    .C(_0615_),
    .D(_1053_),
    .X(_1054_));
 sky130_fd_sc_hd__nor2_1 _2869_ (.A(_0837_),
    .B(_1054_),
    .Y(_1055_));
 sky130_fd_sc_hd__o31a_1 _2870_ (.A1(\usb2uart.u_usb_cdc.endp[0] ),
    .A2(_1047_),
    .A3(_1050_),
    .B1(_1055_),
    .X(_1056_));
 sky130_fd_sc_hd__o31a_1 _2871_ (.A1(\usb2uart.u_usb_cdc.endp[0] ),
    .A2(_1050_),
    .A3(_1046_),
    .B1(_1047_),
    .X(_1057_));
 sky130_fd_sc_hd__o21ba_1 _2872_ (.A1(_1046_),
    .A2(_1056_),
    .B1_N(_1057_),
    .X(_0085_));
 sky130_fd_sc_hd__and2_1 _2873_ (.A(_0518_),
    .B(_0889_),
    .X(_1058_));
 sky130_fd_sc_hd__or3_1 _2874_ (.A(_0597_),
    .B(_0518_),
    .C(\usb2uart.u_usb_cdc.u_sie.phy_state_q[9] ),
    .X(_1059_));
 sky130_fd_sc_hd__or2_2 _2875_ (.A(_2074_),
    .B(_1059_),
    .X(_1060_));
 sky130_fd_sc_hd__a32o_1 _2876_ (.A1(_2003_),
    .A2(_0588_),
    .A3(_1058_),
    .B1(_1060_),
    .B2(\usb2uart.u_usb_cdc.in_data_ack ),
    .X(_0086_));
 sky130_fd_sc_hd__buf_2 _2877_ (.A(_1036_),
    .X(_1061_));
 sky130_fd_sc_hd__nand2_1 _2878_ (.A(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.rx_state_q[2] ),
    .B(_0804_),
    .Y(_1062_));
 sky130_fd_sc_hd__nand2_1 _2879_ (.A(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.rx_state_q[3] ),
    .B(_0810_),
    .Y(_1063_));
 sky130_fd_sc_hd__o31a_1 _2880_ (.A1(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.data_q[0] ),
    .A2(_0821_),
    .A3(_1062_),
    .B1(_1063_),
    .X(_1064_));
 sky130_fd_sc_hd__nor2_2 _2881_ (.A(_1061_),
    .B(_1064_),
    .Y(_1065_));
 sky130_fd_sc_hd__a22o_1 _2882_ (.A1(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.data_q[0] ),
    .A2(_1061_),
    .B1(_1065_),
    .B2(\usb2uart.u_usb_cdc.u_sie.rx_data[0] ),
    .X(_0087_));
 sky130_fd_sc_hd__a22o_1 _2883_ (.A1(\usb2uart.u_usb_cdc.u_sie.rx_data[0] ),
    .A2(_1061_),
    .B1(_1065_),
    .B2(\usb2uart.u_usb_cdc.u_sie.rx_data[1] ),
    .X(_0088_));
 sky130_fd_sc_hd__a22o_1 _2884_ (.A1(\usb2uart.u_usb_cdc.u_sie.rx_data[1] ),
    .A2(_1061_),
    .B1(_1065_),
    .B2(\usb2uart.u_usb_cdc.u_sie.rx_data[2] ),
    .X(_0089_));
 sky130_fd_sc_hd__a22o_1 _2885_ (.A1(\usb2uart.u_usb_cdc.u_sie.rx_data[2] ),
    .A2(_1061_),
    .B1(_1065_),
    .B2(\usb2uart.u_usb_cdc.u_sie.rx_data[3] ),
    .X(_0090_));
 sky130_fd_sc_hd__a22o_1 _2886_ (.A1(\usb2uart.u_usb_cdc.u_sie.rx_data[3] ),
    .A2(_1061_),
    .B1(_1065_),
    .B2(\usb2uart.u_usb_cdc.u_sie.rx_data[4] ),
    .X(_0091_));
 sky130_fd_sc_hd__a22o_1 _2887_ (.A1(\usb2uart.u_usb_cdc.u_sie.rx_data[4] ),
    .A2(_1061_),
    .B1(_1065_),
    .B2(\usb2uart.u_usb_cdc.u_sie.rx_data[5] ),
    .X(_0092_));
 sky130_fd_sc_hd__a22o_1 _2888_ (.A1(\usb2uart.u_usb_cdc.u_sie.rx_data[5] ),
    .A2(_1061_),
    .B1(_1065_),
    .B2(\usb2uart.u_usb_cdc.u_sie.rx_data[6] ),
    .X(_0093_));
 sky130_fd_sc_hd__and3_1 _2889_ (.A(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.rx_state_q[3] ),
    .B(\usb2uart.u_usb_cdc.u_sie.rx_data[7] ),
    .C(_0810_),
    .X(_1066_));
 sky130_fd_sc_hd__o22a_1 _2890_ (.A1(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.data_q[0] ),
    .A2(\usb2uart.u_usb_cdc.u_sie.rx_data[7] ),
    .B1(_1037_),
    .B2(_1066_),
    .X(_1067_));
 sky130_fd_sc_hd__mux2_1 _2891_ (.A0(_1067_),
    .A1(\usb2uart.u_usb_cdc.u_sie.rx_data[6] ),
    .S(_1061_),
    .X(_1068_));
 sky130_fd_sc_hd__clkbuf_1 _2892_ (.A(_1068_),
    .X(_0094_));
 sky130_fd_sc_hd__o211ai_1 _2893_ (.A1(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.rx_state_q[3] ),
    .A2(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.rx_state_q[2] ),
    .B1(_0832_),
    .C1(_1035_),
    .Y(_1069_));
 sky130_fd_sc_hd__mux2_1 _2894_ (.A0(_1069_),
    .A1(\usb2uart.u_usb_cdc.u_sie.rx_data[7] ),
    .S(_1061_),
    .X(_1070_));
 sky130_fd_sc_hd__clkbuf_1 _2895_ (.A(_1070_),
    .X(_0095_));
 sky130_fd_sc_hd__a211o_1 _2896_ (.A1(_0817_),
    .A2(_1062_),
    .B1(_2070_),
    .C1(_0809_),
    .X(_1071_));
 sky130_fd_sc_hd__a21oi_1 _2897_ (.A1(_2065_),
    .A2(_0817_),
    .B1(_1071_),
    .Y(_1072_));
 sky130_fd_sc_hd__mux2_1 _2898_ (.A0(_1072_),
    .A1(_0795_),
    .S(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.stuffing_cnt_q[0] ),
    .X(_1073_));
 sky130_fd_sc_hd__clkbuf_1 _2899_ (.A(_1073_),
    .X(_0096_));
 sky130_fd_sc_hd__nand2_1 _2900_ (.A(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.stuffing_cnt_q[0] ),
    .B(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.stuffing_cnt_q[1] ),
    .Y(_1074_));
 sky130_fd_sc_hd__or2_1 _2901_ (.A(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.stuffing_cnt_q[0] ),
    .B(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.stuffing_cnt_q[1] ),
    .X(_1075_));
 sky130_fd_sc_hd__a32o_1 _2902_ (.A1(_1072_),
    .A2(_1074_),
    .A3(_1075_),
    .B1(_0795_),
    .B2(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.stuffing_cnt_q[1] ),
    .X(_0097_));
 sky130_fd_sc_hd__inv_2 _2903_ (.A(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.stuffing_cnt_q[2] ),
    .Y(_1076_));
 sky130_fd_sc_hd__o211a_1 _2904_ (.A1(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.stuffing_cnt_q[0] ),
    .A2(_0817_),
    .B1(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.stuffing_cnt_q[2] ),
    .C1(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.stuffing_cnt_q[1] ),
    .X(_1077_));
 sky130_fd_sc_hd__o22a_1 _2905_ (.A1(_1076_),
    .A2(_0826_),
    .B1(_1071_),
    .B2(_1077_),
    .X(_1078_));
 sky130_fd_sc_hd__a21oi_1 _2906_ (.A1(_1076_),
    .A2(_1074_),
    .B1(_1078_),
    .Y(_0098_));
 sky130_fd_sc_hd__mux2_1 _2907_ (.A0(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.nrzi_q[2] ),
    .A1(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.nrzi_q[0] ),
    .S(_0795_),
    .X(_1079_));
 sky130_fd_sc_hd__clkbuf_1 _2908_ (.A(_1079_),
    .X(_0099_));
 sky130_fd_sc_hd__mux2_1 _2909_ (.A0(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.nrzi_q[3] ),
    .A1(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.nrzi_q[1] ),
    .S(_0795_),
    .X(_1080_));
 sky130_fd_sc_hd__clkbuf_1 _2910_ (.A(_1080_),
    .X(_0100_));
 sky130_fd_sc_hd__mux2_1 _2911_ (.A0(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.nrzi_q[2] ),
    .A1(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.dp_q[0] ),
    .S(_0826_),
    .X(_1081_));
 sky130_fd_sc_hd__clkbuf_1 _2912_ (.A(_1081_),
    .X(_0101_));
 sky130_fd_sc_hd__mux2_1 _2913_ (.A0(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.nrzi_q[3] ),
    .A1(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.dn_q[0] ),
    .S(_0826_),
    .X(_1082_));
 sky130_fd_sc_hd__clkbuf_1 _2914_ (.A(_1082_),
    .X(_0102_));
 sky130_fd_sc_hd__or4_2 _2915_ (.A(\usb2uart.u_uart.uart_rx_inst.prescale_reg[3] ),
    .B(\usb2uart.u_uart.uart_rx_inst.prescale_reg[2] ),
    .C(\usb2uart.u_uart.uart_rx_inst.prescale_reg[1] ),
    .D(\usb2uart.u_uart.uart_rx_inst.prescale_reg[0] ),
    .X(_1083_));
 sky130_fd_sc_hd__or4_2 _2916_ (.A(\usb2uart.u_uart.uart_rx_inst.prescale_reg[6] ),
    .B(\usb2uart.u_uart.uart_rx_inst.prescale_reg[5] ),
    .C(\usb2uart.u_uart.uart_rx_inst.prescale_reg[4] ),
    .D(_1083_),
    .X(_1084_));
 sky130_fd_sc_hd__or4_2 _2917_ (.A(\usb2uart.u_uart.uart_rx_inst.prescale_reg[9] ),
    .B(\usb2uart.u_uart.uart_rx_inst.prescale_reg[8] ),
    .C(\usb2uart.u_uart.uart_rx_inst.prescale_reg[7] ),
    .D(_1084_),
    .X(_1085_));
 sky130_fd_sc_hd__or4_2 _2918_ (.A(\usb2uart.u_uart.uart_rx_inst.prescale_reg[12] ),
    .B(\usb2uart.u_uart.uart_rx_inst.prescale_reg[11] ),
    .C(\usb2uart.u_uart.uart_rx_inst.prescale_reg[10] ),
    .D(_1085_),
    .X(_1086_));
 sky130_fd_sc_hd__or4_2 _2919_ (.A(\usb2uart.u_uart.uart_rx_inst.prescale_reg[15] ),
    .B(\usb2uart.u_uart.uart_rx_inst.prescale_reg[14] ),
    .C(\usb2uart.u_uart.uart_rx_inst.prescale_reg[13] ),
    .D(_1086_),
    .X(_1087_));
 sky130_fd_sc_hd__or3_1 _2920_ (.A(\usb2uart.u_uart.uart_rx_inst.prescale_reg[17] ),
    .B(\usb2uart.u_uart.uart_rx_inst.prescale_reg[16] ),
    .C(_1087_),
    .X(_1088_));
 sky130_fd_sc_hd__or2_1 _2921_ (.A(\usb2uart.u_uart.uart_rx_inst.prescale_reg[18] ),
    .B(_1088_),
    .X(_1089_));
 sky130_fd_sc_hd__clkbuf_4 _2922_ (.A(_1089_),
    .X(_1090_));
 sky130_fd_sc_hd__nor4_2 _2923_ (.A(\usb2uart.u_uart.uart_rx_inst.bit_cnt[3] ),
    .B(\usb2uart.u_uart.uart_rx_inst.bit_cnt[2] ),
    .C(\usb2uart.u_uart.uart_rx_inst.bit_cnt[1] ),
    .D(_1089_),
    .Y(_1091_));
 sky130_fd_sc_hd__or3_1 _2924_ (.A(\usb2uart.u_uart.uart_rx_inst.bit_cnt[1] ),
    .B(\usb2uart.u_uart.uart_rx_inst.bit_cnt[0] ),
    .C(\usb2uart.u_uart.uart_rx_inst.rxd_reg ),
    .X(_1092_));
 sky130_fd_sc_hd__a21o_2 _2925_ (.A1(_1091_),
    .A2(_1092_),
    .B1(net4),
    .X(_1093_));
 sky130_fd_sc_hd__o21a_1 _2926_ (.A1(\usb2uart.u_uart.uart_rx_inst.bit_cnt[2] ),
    .A2(\usb2uart.u_uart.uart_rx_inst.bit_cnt[1] ),
    .B1(\usb2uart.u_uart.uart_rx_inst.bit_cnt[3] ),
    .X(_1094_));
 sky130_fd_sc_hd__or3_1 _2927_ (.A(_1090_),
    .B(_1093_),
    .C(_1094_),
    .X(_1095_));
 sky130_fd_sc_hd__buf_2 _2928_ (.A(_1095_),
    .X(_1096_));
 sky130_fd_sc_hd__inv_2 _2929_ (.A(\usb2uart.u_uart.uart_rx_inst.bit_cnt[2] ),
    .Y(_1097_));
 sky130_fd_sc_hd__nor2_2 _2930_ (.A(\usb2uart.u_uart.uart_rx_inst.bit_cnt[1] ),
    .B(\usb2uart.u_uart.uart_rx_inst.bit_cnt[0] ),
    .Y(_1098_));
 sky130_fd_sc_hd__and3b_1 _2931_ (.A_N(\usb2uart.u_uart.uart_rx_inst.bit_cnt[3] ),
    .B(_1097_),
    .C(_1098_),
    .X(_1099_));
 sky130_fd_sc_hd__clkbuf_2 _2932_ (.A(_1099_),
    .X(_1100_));
 sky130_fd_sc_hd__nor2_2 _2933_ (.A(_1100_),
    .B(_1096_),
    .Y(_1101_));
 sky130_fd_sc_hd__a22o_1 _2934_ (.A1(\usb2uart.u_uart.uart_rx_inst.data_reg[0] ),
    .A2(_1096_),
    .B1(_1101_),
    .B2(\usb2uart.u_uart.uart_rx_inst.data_reg[1] ),
    .X(_0103_));
 sky130_fd_sc_hd__a22o_1 _2935_ (.A1(\usb2uart.u_uart.uart_rx_inst.data_reg[1] ),
    .A2(_1096_),
    .B1(_1101_),
    .B2(\usb2uart.u_uart.uart_rx_inst.data_reg[2] ),
    .X(_0104_));
 sky130_fd_sc_hd__a22o_1 _2936_ (.A1(\usb2uart.u_uart.uart_rx_inst.data_reg[2] ),
    .A2(_1096_),
    .B1(_1101_),
    .B2(\usb2uart.u_uart.uart_rx_inst.data_reg[3] ),
    .X(_0105_));
 sky130_fd_sc_hd__a22o_1 _2937_ (.A1(\usb2uart.u_uart.uart_rx_inst.data_reg[3] ),
    .A2(_1096_),
    .B1(_1101_),
    .B2(\usb2uart.u_uart.uart_rx_inst.data_reg[4] ),
    .X(_0106_));
 sky130_fd_sc_hd__a22o_1 _2938_ (.A1(\usb2uart.u_uart.uart_rx_inst.data_reg[4] ),
    .A2(_1096_),
    .B1(_1101_),
    .B2(\usb2uart.u_uart.uart_rx_inst.data_reg[5] ),
    .X(_0107_));
 sky130_fd_sc_hd__a22o_1 _2939_ (.A1(\usb2uart.u_uart.uart_rx_inst.data_reg[5] ),
    .A2(_1096_),
    .B1(_1101_),
    .B2(\usb2uart.u_uart.uart_rx_inst.data_reg[6] ),
    .X(_0108_));
 sky130_fd_sc_hd__a22o_1 _2940_ (.A1(\usb2uart.u_uart.uart_rx_inst.data_reg[6] ),
    .A2(_1096_),
    .B1(_1101_),
    .B2(\usb2uart.u_uart.uart_rx_inst.data_reg[7] ),
    .X(_0109_));
 sky130_fd_sc_hd__mux2_1 _2941_ (.A0(\usb2uart.u_uart.uart_rx_inst.rxd_reg ),
    .A1(\usb2uart.u_uart.uart_rx_inst.data_reg[7] ),
    .S(_1096_),
    .X(_1102_));
 sky130_fd_sc_hd__clkbuf_1 _2942_ (.A(_1102_),
    .X(_0110_));
 sky130_fd_sc_hd__or2_1 _2943_ (.A(\usb2uart.u_usb_cdc.u_sie.phy_state_q[8] ),
    .B(_0553_),
    .X(_1103_));
 sky130_fd_sc_hd__o21ai_1 _2944_ (.A1(_0594_),
    .A2(_1103_),
    .B1(_0849_),
    .Y(_1104_));
 sky130_fd_sc_hd__nor2_2 _2945_ (.A(_0553_),
    .B(_0518_),
    .Y(_1105_));
 sky130_fd_sc_hd__o31ai_4 _2946_ (.A1(_0597_),
    .A2(_0633_),
    .A3(_1105_),
    .B1(_0838_),
    .Y(_1106_));
 sky130_fd_sc_hd__mux2_1 _2947_ (.A0(\usb2uart.u_usb_cdc.u_sie.pid_q[0] ),
    .A1(_1104_),
    .S(_1106_),
    .X(_1107_));
 sky130_fd_sc_hd__clkbuf_1 _2948_ (.A(_1107_),
    .X(_0111_));
 sky130_fd_sc_hd__a21o_1 _2949_ (.A1(_0521_),
    .A2(_0527_),
    .B1(_1103_),
    .X(_1108_));
 sky130_fd_sc_hd__mux2_1 _2950_ (.A0(\usb2uart.u_usb_cdc.u_sie.pid_q[1] ),
    .A1(_1108_),
    .S(_1106_),
    .X(_1109_));
 sky130_fd_sc_hd__clkbuf_1 _2951_ (.A(_1109_),
    .X(_0112_));
 sky130_fd_sc_hd__mux2_1 _2952_ (.A0(_0525_),
    .A1(_2055_),
    .S(_1103_),
    .X(_1110_));
 sky130_fd_sc_hd__inv_2 _2953_ (.A(_1110_),
    .Y(_1111_));
 sky130_fd_sc_hd__mux2_1 _2954_ (.A0(\usb2uart.u_usb_cdc.u_sie.pid_q[2] ),
    .A1(_1111_),
    .S(_1106_),
    .X(_1112_));
 sky130_fd_sc_hd__clkbuf_1 _2955_ (.A(_1112_),
    .X(_0113_));
 sky130_fd_sc_hd__inv_2 _2956_ (.A(\usb2uart.u_usb_cdc.bulk_out_nak ),
    .Y(_1113_));
 sky130_fd_sc_hd__o21ai_1 _2957_ (.A1(_1113_),
    .A2(_0861_),
    .B1(_2055_),
    .Y(_1114_));
 sky130_fd_sc_hd__and4b_1 _2958_ (.A_N(\usb2uart.u_usb_cdc.u_sie.phy_state_q[8] ),
    .B(_0630_),
    .C(_0519_),
    .D(_0527_),
    .X(_1115_));
 sky130_fd_sc_hd__a211o_1 _2959_ (.A1(_0553_),
    .A2(_0979_),
    .B1(_1115_),
    .C1(_0631_),
    .X(_1116_));
 sky130_fd_sc_hd__a21o_1 _2960_ (.A1(_0597_),
    .A2(_1114_),
    .B1(_1116_),
    .X(_1117_));
 sky130_fd_sc_hd__mux2_1 _2961_ (.A0(\usb2uart.u_usb_cdc.u_sie.pid_q[3] ),
    .A1(_1117_),
    .S(_1106_),
    .X(_1118_));
 sky130_fd_sc_hd__clkbuf_1 _2962_ (.A(_1118_),
    .X(_0114_));
 sky130_fd_sc_hd__buf_4 _2963_ (.A(_0482_),
    .X(_1119_));
 sky130_fd_sc_hd__or3_1 _2964_ (.A(_2004_),
    .B(_0514_),
    .C(_0576_),
    .X(_1120_));
 sky130_fd_sc_hd__or4_1 _2965_ (.A(_0589_),
    .B(_0593_),
    .C(_1120_),
    .D(_0893_),
    .X(_1121_));
 sky130_fd_sc_hd__buf_4 _2966_ (.A(_1121_),
    .X(_1122_));
 sky130_fd_sc_hd__mux2_1 _2967_ (.A0(_1119_),
    .A1(\usb2uart.u_usb_cdc.u_sie.addr_q[0] ),
    .S(_1122_),
    .X(_1123_));
 sky130_fd_sc_hd__clkbuf_1 _2968_ (.A(_1123_),
    .X(_0115_));
 sky130_fd_sc_hd__clkbuf_4 _2969_ (.A(_0465_),
    .X(_1124_));
 sky130_fd_sc_hd__mux2_1 _2970_ (.A0(_1124_),
    .A1(\usb2uart.u_usb_cdc.u_sie.addr_q[1] ),
    .S(_1122_),
    .X(_1125_));
 sky130_fd_sc_hd__clkbuf_1 _2971_ (.A(_1125_),
    .X(_0116_));
 sky130_fd_sc_hd__buf_4 _2972_ (.A(\usb2uart.u_usb_cdc.out_data[2] ),
    .X(_1126_));
 sky130_fd_sc_hd__mux2_1 _2973_ (.A0(_1126_),
    .A1(\usb2uart.u_usb_cdc.u_sie.addr_q[2] ),
    .S(_1122_),
    .X(_1127_));
 sky130_fd_sc_hd__clkbuf_1 _2974_ (.A(_1127_),
    .X(_0117_));
 sky130_fd_sc_hd__buf_4 _2975_ (.A(\usb2uart.u_usb_cdc.out_data[3] ),
    .X(_1128_));
 sky130_fd_sc_hd__mux2_1 _2976_ (.A0(_1128_),
    .A1(\usb2uart.u_usb_cdc.u_sie.addr_q[3] ),
    .S(_1122_),
    .X(_1129_));
 sky130_fd_sc_hd__clkbuf_1 _2977_ (.A(_1129_),
    .X(_0118_));
 sky130_fd_sc_hd__buf_4 _2978_ (.A(\usb2uart.u_usb_cdc.out_data[4] ),
    .X(_1130_));
 sky130_fd_sc_hd__mux2_1 _2979_ (.A0(_1130_),
    .A1(\usb2uart.u_usb_cdc.u_sie.addr_q[4] ),
    .S(_1122_),
    .X(_1131_));
 sky130_fd_sc_hd__clkbuf_1 _2980_ (.A(_1131_),
    .X(_0119_));
 sky130_fd_sc_hd__clkbuf_4 _2981_ (.A(\usb2uart.u_usb_cdc.out_data[5] ),
    .X(_1132_));
 sky130_fd_sc_hd__mux2_1 _2982_ (.A0(_1132_),
    .A1(\usb2uart.u_usb_cdc.u_sie.addr_q[5] ),
    .S(_1122_),
    .X(_1133_));
 sky130_fd_sc_hd__clkbuf_1 _2983_ (.A(_1133_),
    .X(_0120_));
 sky130_fd_sc_hd__buf_4 _2984_ (.A(_0466_),
    .X(_1134_));
 sky130_fd_sc_hd__mux2_1 _2985_ (.A0(_1134_),
    .A1(\usb2uart.u_usb_cdc.u_sie.addr_q[6] ),
    .S(_1122_),
    .X(_1135_));
 sky130_fd_sc_hd__clkbuf_1 _2986_ (.A(_1135_),
    .X(_0121_));
 sky130_fd_sc_hd__and4b_1 _2987_ (.A_N(_1048_),
    .B(_1113_),
    .C(_0531_),
    .D(_2049_),
    .X(_1136_));
 sky130_fd_sc_hd__a32o_1 _2988_ (.A1(\usb2uart.u_usb_cdc.u_sie.dataout_toggle_q[1] ),
    .A2(\usb2uart.u_usb_cdc.bulk_out_nak ),
    .A3(_2049_),
    .B1(_0516_),
    .B2(_1136_),
    .X(_1137_));
 sky130_fd_sc_hd__or3_1 _2989_ (.A(_0589_),
    .B(_0861_),
    .C(_0837_),
    .X(_1138_));
 sky130_fd_sc_hd__or3b_1 _2990_ (.A(_0736_),
    .B(_0498_),
    .C_N(\usb2uart.u_usb_cdc.in_data_ack ),
    .X(_1139_));
 sky130_fd_sc_hd__or3b_1 _2991_ (.A(_1139_),
    .B(_2019_),
    .C_N(_0643_),
    .X(_1140_));
 sky130_fd_sc_hd__or4_1 _2992_ (.A(_2075_),
    .B(_2006_),
    .C(_0638_),
    .D(_1140_),
    .X(_1141_));
 sky130_fd_sc_hd__and2b_1 _2993_ (.A_N(\usb2uart.u_usb_cdc.u_ctrl_endp.req_q[7] ),
    .B(\usb2uart.u_usb_cdc.u_ctrl_endp.in_endp_q ),
    .X(_1142_));
 sky130_fd_sc_hd__o32a_1 _2994_ (.A1(_1054_),
    .A2(_1050_),
    .A3(_1138_),
    .B1(_1141_),
    .B2(_1142_),
    .X(_1143_));
 sky130_fd_sc_hd__o21a_1 _2995_ (.A1(_0514_),
    .A2(_1143_),
    .B1(\usb2uart.u_usb_cdc.u_sie.dataout_toggle_q[1] ),
    .X(_1144_));
 sky130_fd_sc_hd__a31o_1 _2996_ (.A1(_2003_),
    .A2(_1055_),
    .A3(_1137_),
    .B1(_1144_),
    .X(_0122_));
 sky130_fd_sc_hd__nand2_1 _2997_ (.A(_0844_),
    .B(_0591_),
    .Y(_1145_));
 sky130_fd_sc_hd__buf_2 _2998_ (.A(_0778_),
    .X(_1146_));
 sky130_fd_sc_hd__nand2_2 _2999_ (.A(_0516_),
    .B(_1146_),
    .Y(_1147_));
 sky130_fd_sc_hd__nand2_1 _3000_ (.A(\usb2uart.u_usb_cdc.u_sie.in_byte_q[0] ),
    .B(_1147_),
    .Y(_1148_));
 sky130_fd_sc_hd__o21ai_1 _3001_ (.A1(\usb2uart.u_usb_cdc.u_sie.in_byte_q[0] ),
    .A2(_1145_),
    .B1(_1148_),
    .Y(_0123_));
 sky130_fd_sc_hd__a32o_1 _3002_ (.A1(_0844_),
    .A2(_2053_),
    .A3(_0591_),
    .B1(_1147_),
    .B2(\usb2uart.u_usb_cdc.u_sie.in_byte_q[1] ),
    .X(_1149_));
 sky130_fd_sc_hd__o21a_1 _3003_ (.A1(\usb2uart.u_usb_cdc.u_sie.in_byte_q[1] ),
    .A2(\usb2uart.u_usb_cdc.u_sie.in_byte_q[0] ),
    .B1(_1149_),
    .X(_0124_));
 sky130_fd_sc_hd__o21a_1 _3004_ (.A1(_2052_),
    .A2(_2053_),
    .B1(_0844_),
    .X(_1150_));
 sky130_fd_sc_hd__nor2_1 _3005_ (.A(_2053_),
    .B(_1147_),
    .Y(_1151_));
 sky130_fd_sc_hd__o22a_1 _3006_ (.A1(_1147_),
    .A2(_1150_),
    .B1(_1151_),
    .B2(\usb2uart.u_usb_cdc.u_sie.in_byte_q[2] ),
    .X(_0125_));
 sky130_fd_sc_hd__o21ai_1 _3007_ (.A1(_1147_),
    .A2(_1150_),
    .B1(\usb2uart.u_usb_cdc.u_sie.in_byte_q[3] ),
    .Y(_1152_));
 sky130_fd_sc_hd__o21ai_1 _3008_ (.A1(_2054_),
    .A2(_1145_),
    .B1(_1152_),
    .Y(_0126_));
 sky130_fd_sc_hd__a21oi_1 _3009_ (.A1(\usb2uart.u_usb_cdc.u_sie.delay_cnt_q[0] ),
    .A2(_2074_),
    .B1(_1059_),
    .Y(_0127_));
 sky130_fd_sc_hd__nor3_1 _3010_ (.A(_0597_),
    .B(_0518_),
    .C(\usb2uart.u_usb_cdc.u_sie.phy_state_q[9] ),
    .Y(_1153_));
 sky130_fd_sc_hd__o21ai_1 _3011_ (.A1(\usb2uart.u_usb_cdc.u_sie.delay_cnt_q[1] ),
    .A2(\usb2uart.u_usb_cdc.u_sie.delay_cnt_q[0] ),
    .B1(_1153_),
    .Y(_1154_));
 sky130_fd_sc_hd__a21o_1 _3012_ (.A1(\usb2uart.u_usb_cdc.u_sie.delay_cnt_q[1] ),
    .A2(\usb2uart.u_usb_cdc.u_sie.delay_cnt_q[0] ),
    .B1(_1154_),
    .X(_1155_));
 sky130_fd_sc_hd__nand2_1 _3013_ (.A(_1060_),
    .B(_1155_),
    .Y(_0128_));
 sky130_fd_sc_hd__a21oi_1 _3014_ (.A1(\usb2uart.u_usb_cdc.u_sie.delay_cnt_q[1] ),
    .A2(\usb2uart.u_usb_cdc.u_sie.delay_cnt_q[0] ),
    .B1(\usb2uart.u_usb_cdc.u_sie.delay_cnt_q[2] ),
    .Y(_1156_));
 sky130_fd_sc_hd__o31ai_1 _3015_ (.A1(_2072_),
    .A2(_1059_),
    .A3(_1156_),
    .B1(_1060_),
    .Y(_0129_));
 sky130_fd_sc_hd__inv_2 _3016_ (.A(\usb2uart.u_usb_cdc.u_sie.delay_cnt_q[4] ),
    .Y(_1157_));
 sky130_fd_sc_hd__o21ai_1 _3017_ (.A1(\usb2uart.u_usb_cdc.u_sie.delay_cnt_q[3] ),
    .A2(_2072_),
    .B1(_1153_),
    .Y(_1158_));
 sky130_fd_sc_hd__a21oi_1 _3018_ (.A1(_1157_),
    .A2(_2073_),
    .B1(_1158_),
    .Y(_0130_));
 sky130_fd_sc_hd__o21a_1 _3019_ (.A1(\usb2uart.u_usb_cdc.u_sie.delay_cnt_q[4] ),
    .A2(_2073_),
    .B1(_1153_),
    .X(_0131_));
 sky130_fd_sc_hd__nor2_1 _3020_ (.A(_1054_),
    .B(_1050_),
    .Y(_1159_));
 sky130_fd_sc_hd__a211o_1 _3021_ (.A1(_0597_),
    .A2(_1159_),
    .B1(_1058_),
    .C1(_1044_),
    .X(_1160_));
 sky130_fd_sc_hd__a31o_1 _3022_ (.A1(_2003_),
    .A2(_0588_),
    .A3(_1160_),
    .B1(\usb2uart.u_usb_cdc.u_sie.out_eop_q ),
    .X(_1161_));
 sky130_fd_sc_hd__and2_1 _3023_ (.A(_1060_),
    .B(_1161_),
    .X(_1162_));
 sky130_fd_sc_hd__clkbuf_1 _3024_ (.A(_1162_),
    .X(_0132_));
 sky130_fd_sc_hd__o41a_4 _3025_ (.A1(\usb2uart.u_usb_cdc.u_sie.phy_state_q[7] ),
    .A2(_0553_),
    .A3(_0518_),
    .A4(_0841_),
    .B1(_0590_),
    .X(_1163_));
 sky130_fd_sc_hd__buf_2 _3026_ (.A(_1163_),
    .X(_1164_));
 sky130_fd_sc_hd__nand2_2 _3027_ (.A(_1105_),
    .B(_1163_),
    .Y(_1165_));
 sky130_fd_sc_hd__buf_2 _3028_ (.A(_1165_),
    .X(_1166_));
 sky130_fd_sc_hd__or2_1 _3029_ (.A(_0598_),
    .B(_0612_),
    .X(_1167_));
 sky130_fd_sc_hd__nand2_1 _3030_ (.A(_0613_),
    .B(_1167_),
    .Y(_1168_));
 sky130_fd_sc_hd__o22a_1 _3031_ (.A1(\usb2uart.u_usb_cdc.u_sie.crc16_q[0] ),
    .A2(_1164_),
    .B1(_1166_),
    .B2(_1168_),
    .X(_0133_));
 sky130_fd_sc_hd__o22a_1 _3032_ (.A1(\usb2uart.u_usb_cdc.u_sie.crc16_q[1] ),
    .A2(_1164_),
    .B1(_1166_),
    .B2(_0611_),
    .X(_0134_));
 sky130_fd_sc_hd__o22a_1 _3033_ (.A1(\usb2uart.u_usb_cdc.u_sie.crc16_q[2] ),
    .A2(_1164_),
    .B1(_1166_),
    .B2(_0622_),
    .X(_0135_));
 sky130_fd_sc_hd__o22a_1 _3034_ (.A1(\usb2uart.u_usb_cdc.u_sie.crc16_q[3] ),
    .A2(_1164_),
    .B1(_1166_),
    .B2(_0623_),
    .X(_0136_));
 sky130_fd_sc_hd__o22a_1 _3035_ (.A1(\usb2uart.u_usb_cdc.u_sie.crc16_q[4] ),
    .A2(_1164_),
    .B1(_1166_),
    .B2(_0606_),
    .X(_0137_));
 sky130_fd_sc_hd__o22a_1 _3036_ (.A1(\usb2uart.u_usb_cdc.u_sie.crc16_q[5] ),
    .A2(_1164_),
    .B1(_1166_),
    .B2(_0615_),
    .X(_0138_));
 sky130_fd_sc_hd__o22a_1 _3037_ (.A1(\usb2uart.u_usb_cdc.u_sie.crc16_q[6] ),
    .A2(_1164_),
    .B1(_1166_),
    .B2(_0601_),
    .X(_0139_));
 sky130_fd_sc_hd__o22a_1 _3038_ (.A1(\usb2uart.u_usb_cdc.u_sie.crc16_q[7] ),
    .A2(_1164_),
    .B1(_1166_),
    .B2(_0621_),
    .X(_0140_));
 sky130_fd_sc_hd__o22a_1 _3039_ (.A1(\usb2uart.u_usb_cdc.u_sie.crc16_q[8] ),
    .A2(_1164_),
    .B1(_1166_),
    .B2(_0614_),
    .X(_0141_));
 sky130_fd_sc_hd__o22a_1 _3040_ (.A1(\usb2uart.u_usb_cdc.u_sie.crc16_q[9] ),
    .A2(_1164_),
    .B1(_1166_),
    .B2(_0620_),
    .X(_0142_));
 sky130_fd_sc_hd__o22a_1 _3041_ (.A1(\usb2uart.u_usb_cdc.u_sie.crc16_q[10] ),
    .A2(_1163_),
    .B1(_1165_),
    .B2(\usb2uart.u_usb_cdc.u_sie.crc16_q[2] ),
    .X(_0143_));
 sky130_fd_sc_hd__o22a_1 _3042_ (.A1(\usb2uart.u_usb_cdc.u_sie.crc16_q[11] ),
    .A2(_1163_),
    .B1(_1165_),
    .B2(\usb2uart.u_usb_cdc.u_sie.crc16_q[3] ),
    .X(_0144_));
 sky130_fd_sc_hd__o22a_1 _3043_ (.A1(\usb2uart.u_usb_cdc.u_sie.crc16_q[12] ),
    .A2(_1163_),
    .B1(_1165_),
    .B2(\usb2uart.u_usb_cdc.u_sie.crc16_q[4] ),
    .X(_0145_));
 sky130_fd_sc_hd__o22a_1 _3044_ (.A1(\usb2uart.u_usb_cdc.u_sie.crc16_q[13] ),
    .A2(_1163_),
    .B1(_1165_),
    .B2(\usb2uart.u_usb_cdc.u_sie.crc16_q[5] ),
    .X(_0146_));
 sky130_fd_sc_hd__o22a_1 _3045_ (.A1(\usb2uart.u_usb_cdc.u_sie.crc16_q[14] ),
    .A2(_1163_),
    .B1(_1165_),
    .B2(\usb2uart.u_usb_cdc.u_sie.crc16_q[6] ),
    .X(_0147_));
 sky130_fd_sc_hd__nor2_1 _3046_ (.A(_0955_),
    .B(_1168_),
    .Y(_1169_));
 sky130_fd_sc_hd__and2_1 _3047_ (.A(_0955_),
    .B(_1168_),
    .X(_1170_));
 sky130_fd_sc_hd__o32a_1 _3048_ (.A1(_1165_),
    .A2(_1169_),
    .A3(_1170_),
    .B1(_1163_),
    .B2(\usb2uart.u_usb_cdc.u_sie.crc16_q[15] ),
    .X(_0148_));
 sky130_fd_sc_hd__buf_2 _3049_ (.A(\usb2uart.u_usb_cdc.out_data[7] ),
    .X(_1171_));
 sky130_fd_sc_hd__mux2_1 _3050_ (.A0(_1171_),
    .A1(\usb2uart.u_usb_cdc.endp[0] ),
    .S(_1122_),
    .X(_1172_));
 sky130_fd_sc_hd__clkbuf_1 _3051_ (.A(_1172_),
    .X(_0149_));
 sky130_fd_sc_hd__mux2_1 _3052_ (.A0(_0517_),
    .A1(\usb2uart.u_usb_cdc.endp[1] ),
    .S(_1122_),
    .X(_1173_));
 sky130_fd_sc_hd__clkbuf_1 _3053_ (.A(_1173_),
    .X(_0150_));
 sky130_fd_sc_hd__mux2_1 _3054_ (.A0(_0521_),
    .A1(\usb2uart.u_usb_cdc.endp[2] ),
    .S(_1122_),
    .X(_1174_));
 sky130_fd_sc_hd__clkbuf_1 _3055_ (.A(_1174_),
    .X(_0151_));
 sky130_fd_sc_hd__mux2_1 _3056_ (.A0(\usb2uart.u_usb_cdc.u_sie.data_q[2] ),
    .A1(\usb2uart.u_usb_cdc.endp[3] ),
    .S(_1121_),
    .X(_1175_));
 sky130_fd_sc_hd__clkbuf_1 _3057_ (.A(_1175_),
    .X(_0152_));
 sky130_fd_sc_hd__or4_1 _3058_ (.A(\usb2uart.u_usb_cdc.u_ctrl_endp.addr_q[2] ),
    .B(\usb2uart.u_usb_cdc.u_ctrl_endp.addr_q[5] ),
    .C(\usb2uart.u_usb_cdc.u_ctrl_endp.addr_q[4] ),
    .D(\usb2uart.u_usb_cdc.u_ctrl_endp.addr_q[6] ),
    .X(_1176_));
 sky130_fd_sc_hd__or4_1 _3059_ (.A(\usb2uart.u_usb_cdc.u_ctrl_endp.req_q[7] ),
    .B(\usb2uart.u_usb_cdc.u_ctrl_endp.addr_q[1] ),
    .C(\usb2uart.u_usb_cdc.u_ctrl_endp.addr_q[0] ),
    .D(\usb2uart.u_usb_cdc.u_ctrl_endp.addr_q[3] ),
    .X(_1177_));
 sky130_fd_sc_hd__nor2_1 _3060_ (.A(_1176_),
    .B(_1177_),
    .Y(_1178_));
 sky130_fd_sc_hd__a211o_1 _3061_ (.A1(\usb2uart.u_usb_cdc.u_ctrl_endp.req_q[7] ),
    .A2(\usb2uart.u_usb_cdc.u_ctrl_endp.dev_state_q[0] ),
    .B1(_1178_),
    .C1(\usb2uart.u_usb_cdc.u_ctrl_endp.usb_reset_q ),
    .X(_1179_));
 sky130_fd_sc_hd__o31a_1 _3062_ (.A1(_2017_),
    .A2(_0646_),
    .A3(_0702_),
    .B1(_0473_),
    .X(_1180_));
 sky130_fd_sc_hd__nor3_1 _3063_ (.A(_2081_),
    .B(_0498_),
    .C(_1180_),
    .Y(_1181_));
 sky130_fd_sc_hd__o21a_1 _3064_ (.A1(\usb2uart.u_usb_cdc.u_ctrl_endp.usb_reset_q ),
    .A2(_1181_),
    .B1(_0644_),
    .X(_1182_));
 sky130_fd_sc_hd__mux2_1 _3065_ (.A0(\usb2uart.u_usb_cdc.u_ctrl_endp.dev_state_qq[0] ),
    .A1(_1179_),
    .S(_1182_),
    .X(_1183_));
 sky130_fd_sc_hd__clkbuf_1 _3066_ (.A(_1183_),
    .X(_0153_));
 sky130_fd_sc_hd__inv_2 _3067_ (.A(\usb2uart.u_usb_cdc.u_ctrl_endp.dev_state_q[1] ),
    .Y(_1184_));
 sky130_fd_sc_hd__a211oi_1 _3068_ (.A1(\usb2uart.u_usb_cdc.u_ctrl_endp.req_q[7] ),
    .A2(_1184_),
    .B1(_1178_),
    .C1(\usb2uart.u_usb_cdc.u_ctrl_endp.usb_reset_q ),
    .Y(_1185_));
 sky130_fd_sc_hd__mux2_1 _3069_ (.A0(\usb2uart.u_usb_cdc.u_ctrl_endp.dev_state_qq[1] ),
    .A1(_1185_),
    .S(_1182_),
    .X(_1186_));
 sky130_fd_sc_hd__clkbuf_1 _3070_ (.A(_1186_),
    .X(_0154_));
 sky130_fd_sc_hd__o21ai_1 _3071_ (.A1(_2004_),
    .A2(_1159_),
    .B1(_2003_),
    .Y(_1187_));
 sky130_fd_sc_hd__a22o_1 _3072_ (.A1(_0652_),
    .A2(_1060_),
    .B1(_1187_),
    .B2(_0597_),
    .X(_0155_));
 sky130_fd_sc_hd__buf_2 _3073_ (.A(_2023_),
    .X(_1188_));
 sky130_fd_sc_hd__buf_2 _3074_ (.A(_1188_),
    .X(_1189_));
 sky130_fd_sc_hd__nand2_1 _3075_ (.A(_0452_),
    .B(_0700_),
    .Y(_1190_));
 sky130_fd_sc_hd__clkinv_2 _3076_ (.A(\usb2uart.u_usb_cdc.u_ctrl_endp.req_q[8] ),
    .Y(_1191_));
 sky130_fd_sc_hd__nor2_2 _3077_ (.A(_0452_),
    .B(_1191_),
    .Y(_1192_));
 sky130_fd_sc_hd__o21ai_1 _3078_ (.A1(_0492_),
    .A2(_0480_),
    .B1(_1192_),
    .Y(_1193_));
 sky130_fd_sc_hd__o21a_1 _3079_ (.A1(_2083_),
    .A2(_1190_),
    .B1(_1193_),
    .X(_1194_));
 sky130_fd_sc_hd__nor2_1 _3080_ (.A(_1191_),
    .B(_0478_),
    .Y(_1195_));
 sky130_fd_sc_hd__nand2_1 _3081_ (.A(_0452_),
    .B(_1195_),
    .Y(_1196_));
 sky130_fd_sc_hd__or2_1 _3082_ (.A(_0453_),
    .B(_1196_),
    .X(_1197_));
 sky130_fd_sc_hd__a21oi_1 _3083_ (.A1(_1194_),
    .A2(_1197_),
    .B1(_2026_),
    .Y(_1198_));
 sky130_fd_sc_hd__mux2_1 _3084_ (.A0(_0492_),
    .A1(_0480_),
    .S(_0453_),
    .X(_1199_));
 sky130_fd_sc_hd__nand2_1 _3085_ (.A(_1188_),
    .B(_1199_),
    .Y(_1200_));
 sky130_fd_sc_hd__a21oi_1 _3086_ (.A1(_1188_),
    .A2(_1190_),
    .B1(_2024_),
    .Y(_1201_));
 sky130_fd_sc_hd__o211a_1 _3087_ (.A1(_1189_),
    .A2(_1198_),
    .B1(_1200_),
    .C1(_1201_),
    .X(_1202_));
 sky130_fd_sc_hd__or3_1 _3088_ (.A(_2084_),
    .B(_0450_),
    .C(_0760_),
    .X(_1203_));
 sky130_fd_sc_hd__o211a_1 _3089_ (.A1(_2083_),
    .A2(_1191_),
    .B1(_2040_),
    .C1(_1203_),
    .X(_1204_));
 sky130_fd_sc_hd__buf_2 _3090_ (.A(_0452_),
    .X(_1205_));
 sky130_fd_sc_hd__nand2_1 _3091_ (.A(_0700_),
    .B(_0451_),
    .Y(_1206_));
 sky130_fd_sc_hd__o311a_1 _3092_ (.A1(_2084_),
    .A2(_0452_),
    .A3(_0700_),
    .B1(_0478_),
    .C1(_0453_),
    .X(_1207_));
 sky130_fd_sc_hd__a31o_1 _3093_ (.A1(_1205_),
    .A2(_0639_),
    .A3(_1206_),
    .B1(_1207_),
    .X(_1208_));
 sky130_fd_sc_hd__buf_2 _3094_ (.A(_0453_),
    .X(_1209_));
 sky130_fd_sc_hd__nand2_1 _3095_ (.A(_2083_),
    .B(_1192_),
    .Y(_1210_));
 sky130_fd_sc_hd__nand2_1 _3096_ (.A(_0450_),
    .B(_0700_),
    .Y(_1211_));
 sky130_fd_sc_hd__a22o_1 _3097_ (.A1(_1209_),
    .A2(_1210_),
    .B1(_1211_),
    .B2(_1205_),
    .X(_1212_));
 sky130_fd_sc_hd__mux2_1 _3098_ (.A0(_1208_),
    .A1(_1212_),
    .S(_1188_),
    .X(_1213_));
 sky130_fd_sc_hd__nor3_1 _3099_ (.A(_0454_),
    .B(_1204_),
    .C(_1213_),
    .Y(_1214_));
 sky130_fd_sc_hd__or4b_1 _3100_ (.A(_2006_),
    .B(_0883_),
    .C(_2081_),
    .D_N(\usb2uart.u_usb_cdc.u_ctrl_endp.state_q[3] ),
    .X(_1215_));
 sky130_fd_sc_hd__nor2_1 _3101_ (.A(_0655_),
    .B(_1215_),
    .Y(_1216_));
 sky130_fd_sc_hd__and3b_2 _3102_ (.A_N(\usb2uart.u_usb_cdc.u_ctrl_endp.byte_cnt_q[6] ),
    .B(_0701_),
    .C(_1216_),
    .X(_1217_));
 sky130_fd_sc_hd__o21a_1 _3103_ (.A1(_1202_),
    .A2(_1214_),
    .B1(_1217_),
    .X(_1218_));
 sky130_fd_sc_hd__inv_2 _3104_ (.A(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_first_qq[3] ),
    .Y(_1219_));
 sky130_fd_sc_hd__buf_2 _3105_ (.A(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_first_qq[1] ),
    .X(_1220_));
 sky130_fd_sc_hd__buf_2 _3106_ (.A(_1220_),
    .X(_1221_));
 sky130_fd_sc_hd__buf_4 _3107_ (.A(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_first_qq[0] ),
    .X(_1222_));
 sky130_fd_sc_hd__buf_4 _3108_ (.A(_1222_),
    .X(_1223_));
 sky130_fd_sc_hd__mux2_1 _3109_ (.A0(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[48] ),
    .A1(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[56] ),
    .S(_1223_),
    .X(_1224_));
 sky130_fd_sc_hd__mux2_1 _3110_ (.A0(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[32] ),
    .A1(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[40] ),
    .S(_1222_),
    .X(_1225_));
 sky130_fd_sc_hd__inv_2 _3111_ (.A(_1225_),
    .Y(_1226_));
 sky130_fd_sc_hd__buf_2 _3112_ (.A(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_first_qq[2] ),
    .X(_1227_));
 sky130_fd_sc_hd__o21ai_1 _3113_ (.A1(_1220_),
    .A2(_1226_),
    .B1(_1227_),
    .Y(_1228_));
 sky130_fd_sc_hd__a21o_1 _3114_ (.A1(_1221_),
    .A2(_1224_),
    .B1(_1228_),
    .X(_1229_));
 sky130_fd_sc_hd__mux2_1 _3115_ (.A0(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[16] ),
    .A1(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[24] ),
    .S(_1223_),
    .X(_1230_));
 sky130_fd_sc_hd__mux2_1 _3116_ (.A0(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[0] ),
    .A1(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[8] ),
    .S(_1222_),
    .X(_1231_));
 sky130_fd_sc_hd__and2b_1 _3117_ (.A_N(_1220_),
    .B(_1231_),
    .X(_1232_));
 sky130_fd_sc_hd__a211o_1 _3118_ (.A1(_1220_),
    .A2(_1230_),
    .B1(_1232_),
    .C1(_1227_),
    .X(_1233_));
 sky130_fd_sc_hd__nor2_1 _3119_ (.A(_1222_),
    .B(_1220_),
    .Y(_1234_));
 sky130_fd_sc_hd__and3b_2 _3120_ (.A_N(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_first_qq[2] ),
    .B(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_first_qq[3] ),
    .C(_1234_),
    .X(_1235_));
 sky130_fd_sc_hd__a32o_1 _3121_ (.A1(_1219_),
    .A2(_1229_),
    .A3(_1233_),
    .B1(_1235_),
    .B2(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[64] ),
    .X(_1236_));
 sky130_fd_sc_hd__a32o_1 _3122_ (.A1(\usb2uart.u_usb_cdc.u_ctrl_endp.req_q[3] ),
    .A2(_0709_),
    .A3(_1216_),
    .B1(_1236_),
    .B2(_0883_),
    .X(_1237_));
 sky130_fd_sc_hd__or3_1 _3123_ (.A(_0884_),
    .B(_1218_),
    .C(_1237_),
    .X(_1238_));
 sky130_fd_sc_hd__o21a_1 _3124_ (.A1(\usb2uart.u_usb_cdc.u_sie.rx_data[0] ),
    .A2(_1146_),
    .B1(_0836_),
    .X(_1239_));
 sky130_fd_sc_hd__a22o_1 _3125_ (.A1(_0517_),
    .A2(_0515_),
    .B1(_1238_),
    .B2(_1239_),
    .X(_0156_));
 sky130_fd_sc_hd__buf_2 _3126_ (.A(_1209_),
    .X(_1240_));
 sky130_fd_sc_hd__nor2_1 _3127_ (.A(_1205_),
    .B(_0480_),
    .Y(_1241_));
 sky130_fd_sc_hd__nand2_1 _3128_ (.A(_2083_),
    .B(_0450_),
    .Y(_1242_));
 sky130_fd_sc_hd__a21oi_1 _3129_ (.A1(_0641_),
    .A2(_1242_),
    .B1(_0700_),
    .Y(_1243_));
 sky130_fd_sc_hd__and2b_1 _3130_ (.A_N(_0452_),
    .B(_1243_),
    .X(_1244_));
 sky130_fd_sc_hd__a311o_1 _3131_ (.A1(_0760_),
    .A2(_0641_),
    .A3(_1241_),
    .B1(_1244_),
    .C1(_0493_),
    .X(_1245_));
 sky130_fd_sc_hd__nor2_1 _3132_ (.A(_1191_),
    .B(_0641_),
    .Y(_1246_));
 sky130_fd_sc_hd__nor2_1 _3133_ (.A(_0452_),
    .B(_1246_),
    .Y(_1247_));
 sky130_fd_sc_hd__a21o_1 _3134_ (.A1(_1205_),
    .A2(_1211_),
    .B1(_1247_),
    .X(_1248_));
 sky130_fd_sc_hd__o41a_1 _3135_ (.A1(_2083_),
    .A2(_0477_),
    .A3(_0639_),
    .A4(_1190_),
    .B1(_1188_),
    .X(_1249_));
 sky130_fd_sc_hd__a21oi_1 _3136_ (.A1(_1240_),
    .A2(_1248_),
    .B1(_1249_),
    .Y(_1250_));
 sky130_fd_sc_hd__o21a_1 _3137_ (.A1(_1240_),
    .A2(_1245_),
    .B1(_1250_),
    .X(_1251_));
 sky130_fd_sc_hd__a21oi_1 _3138_ (.A1(_1205_),
    .A2(_1206_),
    .B1(_1209_),
    .Y(_1252_));
 sky130_fd_sc_hd__o211a_1 _3139_ (.A1(_0492_),
    .A2(_0502_),
    .B1(_0453_),
    .C1(_0700_),
    .X(_1253_));
 sky130_fd_sc_hd__a31o_1 _3140_ (.A1(_0477_),
    .A2(_0760_),
    .A3(_1252_),
    .B1(_1253_),
    .X(_1254_));
 sky130_fd_sc_hd__a21o_1 _3141_ (.A1(_2039_),
    .A2(_1192_),
    .B1(_0453_),
    .X(_1255_));
 sky130_fd_sc_hd__a31o_1 _3142_ (.A1(_2083_),
    .A2(_1205_),
    .A3(_0760_),
    .B1(_1255_),
    .X(_1256_));
 sky130_fd_sc_hd__a21oi_1 _3143_ (.A1(_1209_),
    .A2(_1193_),
    .B1(_1188_),
    .Y(_1257_));
 sky130_fd_sc_hd__a221o_1 _3144_ (.A1(_1189_),
    .A2(_1254_),
    .B1(_1256_),
    .B2(_1257_),
    .C1(_2024_),
    .X(_1258_));
 sky130_fd_sc_hd__o21a_1 _3145_ (.A1(_0454_),
    .A2(_1251_),
    .B1(_1258_),
    .X(_1259_));
 sky130_fd_sc_hd__clkbuf_4 _3146_ (.A(_1221_),
    .X(_1260_));
 sky130_fd_sc_hd__buf_4 _3147_ (.A(_1222_),
    .X(_1261_));
 sky130_fd_sc_hd__mux2_1 _3148_ (.A0(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[17] ),
    .A1(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[25] ),
    .S(_1261_),
    .X(_1262_));
 sky130_fd_sc_hd__mux2_1 _3149_ (.A0(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[1] ),
    .A1(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[9] ),
    .S(_1223_),
    .X(_1263_));
 sky130_fd_sc_hd__and2b_1 _3150_ (.A_N(_1221_),
    .B(_1263_),
    .X(_1264_));
 sky130_fd_sc_hd__clkbuf_4 _3151_ (.A(_1227_),
    .X(_1265_));
 sky130_fd_sc_hd__a211o_1 _3152_ (.A1(_1260_),
    .A2(_1262_),
    .B1(_1264_),
    .C1(_1265_),
    .X(_1266_));
 sky130_fd_sc_hd__buf_2 _3153_ (.A(_1261_),
    .X(_1267_));
 sky130_fd_sc_hd__mux2_1 _3154_ (.A0(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[49] ),
    .A1(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[57] ),
    .S(_1267_),
    .X(_1268_));
 sky130_fd_sc_hd__buf_2 _3155_ (.A(_1220_),
    .X(_1269_));
 sky130_fd_sc_hd__mux2_1 _3156_ (.A0(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[33] ),
    .A1(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[41] ),
    .S(_1222_),
    .X(_1270_));
 sky130_fd_sc_hd__inv_2 _3157_ (.A(_1270_),
    .Y(_1271_));
 sky130_fd_sc_hd__o21ai_1 _3158_ (.A1(_1269_),
    .A2(_1271_),
    .B1(_1227_),
    .Y(_1272_));
 sky130_fd_sc_hd__a21o_1 _3159_ (.A1(_1260_),
    .A2(_1268_),
    .B1(_1272_),
    .X(_1273_));
 sky130_fd_sc_hd__a32o_1 _3160_ (.A1(_1219_),
    .A2(_1266_),
    .A3(_1273_),
    .B1(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[65] ),
    .B2(_1235_),
    .X(_1274_));
 sky130_fd_sc_hd__a221o_1 _3161_ (.A1(_1217_),
    .A2(_1259_),
    .B1(_1274_),
    .B2(_0883_),
    .C1(_0884_),
    .X(_1275_));
 sky130_fd_sc_hd__o21a_1 _3162_ (.A1(\usb2uart.u_usb_cdc.u_sie.rx_data[1] ),
    .A2(_1146_),
    .B1(_0836_),
    .X(_1276_));
 sky130_fd_sc_hd__a22o_1 _3163_ (.A1(_0521_),
    .A2(_0515_),
    .B1(_1275_),
    .B2(_1276_),
    .X(_0157_));
 sky130_fd_sc_hd__a21oi_1 _3164_ (.A1(_2025_),
    .A2(_1196_),
    .B1(_1188_),
    .Y(_1277_));
 sky130_fd_sc_hd__a211o_1 _3165_ (.A1(_0477_),
    .A2(_1189_),
    .B1(_1277_),
    .C1(_0639_),
    .X(_1278_));
 sky130_fd_sc_hd__a31o_1 _3166_ (.A1(_0760_),
    .A2(_1242_),
    .A3(_0494_),
    .B1(_1240_),
    .X(_1279_));
 sky130_fd_sc_hd__o31ai_1 _3167_ (.A1(_0450_),
    .A2(_1191_),
    .A3(_1247_),
    .B1(_1209_),
    .Y(_1280_));
 sky130_fd_sc_hd__a21o_1 _3168_ (.A1(_0760_),
    .A2(_0502_),
    .B1(_0453_),
    .X(_1281_));
 sky130_fd_sc_hd__a21o_1 _3169_ (.A1(_0450_),
    .A2(_1192_),
    .B1(_1281_),
    .X(_1282_));
 sky130_fd_sc_hd__o21ai_1 _3170_ (.A1(_2084_),
    .A2(_0760_),
    .B1(_1211_),
    .Y(_1283_));
 sky130_fd_sc_hd__and4b_1 _3171_ (.A_N(_1188_),
    .B(_1241_),
    .C(_1283_),
    .D(_1209_),
    .X(_1284_));
 sky130_fd_sc_hd__a31o_1 _3172_ (.A1(_1189_),
    .A2(_1280_),
    .A3(_1282_),
    .B1(_1284_),
    .X(_1285_));
 sky130_fd_sc_hd__a32o_1 _3173_ (.A1(_1201_),
    .A2(_1278_),
    .A3(_1279_),
    .B1(_1285_),
    .B2(_2024_),
    .X(_1286_));
 sky130_fd_sc_hd__mux2_1 _3174_ (.A0(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[18] ),
    .A1(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[26] ),
    .S(_1261_),
    .X(_1287_));
 sky130_fd_sc_hd__mux2_1 _3175_ (.A0(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[2] ),
    .A1(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[10] ),
    .S(_1223_),
    .X(_1288_));
 sky130_fd_sc_hd__and2b_1 _3176_ (.A_N(_1221_),
    .B(_1288_),
    .X(_1289_));
 sky130_fd_sc_hd__a211o_1 _3177_ (.A1(_1260_),
    .A2(_1287_),
    .B1(_1289_),
    .C1(_1265_),
    .X(_1290_));
 sky130_fd_sc_hd__mux2_1 _3178_ (.A0(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[50] ),
    .A1(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[58] ),
    .S(_1267_),
    .X(_1291_));
 sky130_fd_sc_hd__mux2_1 _3179_ (.A0(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[34] ),
    .A1(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[42] ),
    .S(_1222_),
    .X(_1292_));
 sky130_fd_sc_hd__inv_2 _3180_ (.A(_1292_),
    .Y(_1293_));
 sky130_fd_sc_hd__o21ai_1 _3181_ (.A1(_1269_),
    .A2(_1293_),
    .B1(_1227_),
    .Y(_1294_));
 sky130_fd_sc_hd__a21o_1 _3182_ (.A1(_1260_),
    .A2(_1291_),
    .B1(_1294_),
    .X(_1295_));
 sky130_fd_sc_hd__a32o_1 _3183_ (.A1(_1219_),
    .A2(_1290_),
    .A3(_1295_),
    .B1(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[66] ),
    .B2(_1235_),
    .X(_1296_));
 sky130_fd_sc_hd__a221o_1 _3184_ (.A1(_1217_),
    .A2(_1286_),
    .B1(_1296_),
    .B2(_0883_),
    .C1(_0884_),
    .X(_1297_));
 sky130_fd_sc_hd__o21a_1 _3185_ (.A1(\usb2uart.u_usb_cdc.u_sie.rx_data[2] ),
    .A2(_1146_),
    .B1(_0836_),
    .X(_1298_));
 sky130_fd_sc_hd__a22o_1 _3186_ (.A1(\usb2uart.u_usb_cdc.u_sie.data_q[2] ),
    .A2(_0515_),
    .B1(_1297_),
    .B2(_1298_),
    .X(_0158_));
 sky130_fd_sc_hd__mux2_1 _3187_ (.A0(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[35] ),
    .A1(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[43] ),
    .S(_1223_),
    .X(_1299_));
 sky130_fd_sc_hd__or2b_1 _3188_ (.A(_1221_),
    .B_N(_1299_),
    .X(_1300_));
 sky130_fd_sc_hd__mux2_1 _3189_ (.A0(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[51] ),
    .A1(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[59] ),
    .S(_1261_),
    .X(_1301_));
 sky130_fd_sc_hd__nand2_1 _3190_ (.A(_1269_),
    .B(_1301_),
    .Y(_1302_));
 sky130_fd_sc_hd__mux2_1 _3191_ (.A0(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[3] ),
    .A1(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[11] ),
    .S(_1261_),
    .X(_1303_));
 sky130_fd_sc_hd__or2b_1 _3192_ (.A(_1221_),
    .B_N(_1303_),
    .X(_1304_));
 sky130_fd_sc_hd__mux2_1 _3193_ (.A0(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[19] ),
    .A1(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[27] ),
    .S(_1261_),
    .X(_1305_));
 sky130_fd_sc_hd__a21oi_1 _3194_ (.A1(_1269_),
    .A2(_1305_),
    .B1(_1227_),
    .Y(_1306_));
 sky130_fd_sc_hd__a32o_1 _3195_ (.A1(_1265_),
    .A2(_1300_),
    .A3(_1302_),
    .B1(_1304_),
    .B2(_1306_),
    .X(_1307_));
 sky130_fd_sc_hd__o2bb2a_1 _3196_ (.A1_N(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[67] ),
    .A2_N(_1235_),
    .B1(_1307_),
    .B2(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_first_qq[3] ),
    .X(_1308_));
 sky130_fd_sc_hd__nor2_2 _3197_ (.A(\usb2uart.u_usb_cdc.u_ctrl_endp.req_q[2] ),
    .B(_0760_),
    .Y(_1309_));
 sky130_fd_sc_hd__nand2_1 _3198_ (.A(_0700_),
    .B(_0493_),
    .Y(_1310_));
 sky130_fd_sc_hd__a211oi_1 _3199_ (.A1(_1210_),
    .A2(_1310_),
    .B1(_0639_),
    .C1(_2023_),
    .Y(_1311_));
 sky130_fd_sc_hd__a31o_1 _3200_ (.A1(_2023_),
    .A2(_1192_),
    .A3(_0451_),
    .B1(_1311_),
    .X(_1312_));
 sky130_fd_sc_hd__nand2_1 _3201_ (.A(_0454_),
    .B(_1312_),
    .Y(_1313_));
 sky130_fd_sc_hd__a2bb2o_1 _3202_ (.A1_N(_1192_),
    .A2_N(_0502_),
    .B1(_0700_),
    .B2(_0641_),
    .X(_1314_));
 sky130_fd_sc_hd__or4_1 _3203_ (.A(_1209_),
    .B(_2023_),
    .C(_0454_),
    .D(_1314_),
    .X(_1315_));
 sky130_fd_sc_hd__o211a_1 _3204_ (.A1(_2015_),
    .A2(_0478_),
    .B1(_1313_),
    .C1(_1315_),
    .X(_1316_));
 sky130_fd_sc_hd__o31a_1 _3205_ (.A1(_1205_),
    .A2(_1209_),
    .A3(_0641_),
    .B1(\usb2uart.u_usb_cdc.u_ctrl_endp.byte_cnt_q[6] ),
    .X(_1317_));
 sky130_fd_sc_hd__or4b_1 _3206_ (.A(_1309_),
    .B(_1316_),
    .C(_1317_),
    .D_N(_1216_),
    .X(_1318_));
 sky130_fd_sc_hd__o211a_1 _3207_ (.A1(_2009_),
    .A2(_1308_),
    .B1(_1318_),
    .C1(_1146_),
    .X(_1319_));
 sky130_fd_sc_hd__o21ai_1 _3208_ (.A1(\usb2uart.u_usb_cdc.u_sie.rx_data[3] ),
    .A2(_1146_),
    .B1(_0836_),
    .Y(_1320_));
 sky130_fd_sc_hd__a2bb2o_1 _3209_ (.A1_N(_1319_),
    .A2_N(_1320_),
    .B1(_0519_),
    .B2(_0515_),
    .X(_0159_));
 sky130_fd_sc_hd__mux2_1 _3210_ (.A0(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[20] ),
    .A1(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[28] ),
    .S(_1261_),
    .X(_1321_));
 sky130_fd_sc_hd__mux2_1 _3211_ (.A0(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[4] ),
    .A1(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[12] ),
    .S(_1223_),
    .X(_1322_));
 sky130_fd_sc_hd__and2b_1 _3212_ (.A_N(_1221_),
    .B(_1322_),
    .X(_1323_));
 sky130_fd_sc_hd__a211o_1 _3213_ (.A1(_1260_),
    .A2(_1321_),
    .B1(_1323_),
    .C1(_1265_),
    .X(_1324_));
 sky130_fd_sc_hd__mux2_1 _3214_ (.A0(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[52] ),
    .A1(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[60] ),
    .S(_1267_),
    .X(_1325_));
 sky130_fd_sc_hd__mux2_1 _3215_ (.A0(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[36] ),
    .A1(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[44] ),
    .S(_1223_),
    .X(_1326_));
 sky130_fd_sc_hd__inv_2 _3216_ (.A(_1326_),
    .Y(_1327_));
 sky130_fd_sc_hd__o21ai_1 _3217_ (.A1(_1269_),
    .A2(_1327_),
    .B1(_1227_),
    .Y(_1328_));
 sky130_fd_sc_hd__a21o_1 _3218_ (.A1(_1260_),
    .A2(_1325_),
    .B1(_1328_),
    .X(_1329_));
 sky130_fd_sc_hd__a32o_1 _3219_ (.A1(_1219_),
    .A2(_1324_),
    .A3(_1329_),
    .B1(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[68] ),
    .B2(_1235_),
    .X(_1330_));
 sky130_fd_sc_hd__a21oi_1 _3220_ (.A1(_0760_),
    .A2(_0641_),
    .B1(_1189_),
    .Y(_1331_));
 sky130_fd_sc_hd__o211a_1 _3221_ (.A1(_1240_),
    .A2(_1243_),
    .B1(_1241_),
    .C1(_1331_),
    .X(_1332_));
 sky130_fd_sc_hd__a41o_1 _3222_ (.A1(_1205_),
    .A2(_0639_),
    .A3(_1189_),
    .A4(_1195_),
    .B1(_0454_),
    .X(_1333_));
 sky130_fd_sc_hd__o31ai_1 _3223_ (.A1(_0639_),
    .A2(_1188_),
    .A3(_2025_),
    .B1(_0454_),
    .Y(_1334_));
 sky130_fd_sc_hd__o211a_1 _3224_ (.A1(_1332_),
    .A2(_1333_),
    .B1(_1334_),
    .C1(_1217_),
    .X(_1335_));
 sky130_fd_sc_hd__a211o_1 _3225_ (.A1(_0883_),
    .A2(_1330_),
    .B1(_1335_),
    .C1(_0884_),
    .X(_1336_));
 sky130_fd_sc_hd__o21a_1 _3226_ (.A1(\usb2uart.u_usb_cdc.u_sie.rx_data[4] ),
    .A2(_1146_),
    .B1(_0836_),
    .X(_1337_));
 sky130_fd_sc_hd__a22o_1 _3227_ (.A1(\usb2uart.u_usb_cdc.u_sie.data_q[4] ),
    .A2(_0515_),
    .B1(_1336_),
    .B2(_1337_),
    .X(_0160_));
 sky130_fd_sc_hd__a21oi_1 _3228_ (.A1(_1205_),
    .A2(_1206_),
    .B1(_1247_),
    .Y(_1338_));
 sky130_fd_sc_hd__a21o_1 _3229_ (.A1(_1240_),
    .A2(_1338_),
    .B1(_2026_),
    .X(_1339_));
 sky130_fd_sc_hd__a21oi_1 _3230_ (.A1(_0450_),
    .A2(_1191_),
    .B1(_1246_),
    .Y(_1340_));
 sky130_fd_sc_hd__a21oi_1 _3231_ (.A1(_1192_),
    .A2(_0451_),
    .B1(_1209_),
    .Y(_1341_));
 sky130_fd_sc_hd__nand2_1 _3232_ (.A(_1209_),
    .B(_2025_),
    .Y(_1342_));
 sky130_fd_sc_hd__or4b_1 _3233_ (.A(_1188_),
    .B(_2024_),
    .C(_1341_),
    .D_N(_1342_),
    .X(_1343_));
 sky130_fd_sc_hd__o21ai_1 _3234_ (.A1(_2015_),
    .A2(_1340_),
    .B1(_1343_),
    .Y(_1344_));
 sky130_fd_sc_hd__a31o_1 _3235_ (.A1(_1189_),
    .A2(_2024_),
    .A3(_1339_),
    .B1(_1344_),
    .X(_1345_));
 sky130_fd_sc_hd__mux2_1 _3236_ (.A0(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[21] ),
    .A1(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[29] ),
    .S(_1261_),
    .X(_1346_));
 sky130_fd_sc_hd__mux2_1 _3237_ (.A0(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[5] ),
    .A1(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[13] ),
    .S(_1223_),
    .X(_1347_));
 sky130_fd_sc_hd__and2b_1 _3238_ (.A_N(_1221_),
    .B(_1347_),
    .X(_1348_));
 sky130_fd_sc_hd__a211o_1 _3239_ (.A1(_1269_),
    .A2(_1346_),
    .B1(_1348_),
    .C1(_1265_),
    .X(_1349_));
 sky130_fd_sc_hd__mux2_1 _3240_ (.A0(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[53] ),
    .A1(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[61] ),
    .S(_1267_),
    .X(_1350_));
 sky130_fd_sc_hd__mux2_1 _3241_ (.A0(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[37] ),
    .A1(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[45] ),
    .S(_1222_),
    .X(_1351_));
 sky130_fd_sc_hd__inv_2 _3242_ (.A(_1351_),
    .Y(_1352_));
 sky130_fd_sc_hd__o21ai_1 _3243_ (.A1(_1269_),
    .A2(_1352_),
    .B1(_1227_),
    .Y(_1353_));
 sky130_fd_sc_hd__a21o_1 _3244_ (.A1(_1260_),
    .A2(_1350_),
    .B1(_1353_),
    .X(_1354_));
 sky130_fd_sc_hd__a32o_1 _3245_ (.A1(_1219_),
    .A2(_1349_),
    .A3(_1354_),
    .B1(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[69] ),
    .B2(_1235_),
    .X(_1355_));
 sky130_fd_sc_hd__a221o_1 _3246_ (.A1(_1217_),
    .A2(_1345_),
    .B1(_1355_),
    .B2(_0883_),
    .C1(_0884_),
    .X(_1356_));
 sky130_fd_sc_hd__o21a_1 _3247_ (.A1(\usb2uart.u_usb_cdc.u_sie.rx_data[5] ),
    .A2(_1146_),
    .B1(_0836_),
    .X(_1357_));
 sky130_fd_sc_hd__a22o_1 _3248_ (.A1(\usb2uart.u_usb_cdc.u_sie.data_q[5] ),
    .A2(_0515_),
    .B1(_1356_),
    .B2(_1357_),
    .X(_0161_));
 sky130_fd_sc_hd__o21ba_1 _3249_ (.A1(_0639_),
    .A2(_1244_),
    .B1_N(_2023_),
    .X(_1358_));
 sky130_fd_sc_hd__a21o_1 _3250_ (.A1(_1255_),
    .A2(_1358_),
    .B1(_0454_),
    .X(_1359_));
 sky130_fd_sc_hd__mux2_1 _3251_ (.A0(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[38] ),
    .A1(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[46] ),
    .S(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_first_qq[0] ),
    .X(_1360_));
 sky130_fd_sc_hd__or2b_1 _3252_ (.A(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_first_qq[1] ),
    .B_N(_1360_),
    .X(_1361_));
 sky130_fd_sc_hd__mux2_1 _3253_ (.A0(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[54] ),
    .A1(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[62] ),
    .S(_1222_),
    .X(_1362_));
 sky130_fd_sc_hd__nand2_1 _3254_ (.A(_1220_),
    .B(_1362_),
    .Y(_1363_));
 sky130_fd_sc_hd__mux2_1 _3255_ (.A0(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[6] ),
    .A1(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[14] ),
    .S(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_first_qq[0] ),
    .X(_1364_));
 sky130_fd_sc_hd__or2b_1 _3256_ (.A(_1220_),
    .B_N(_1364_),
    .X(_1365_));
 sky130_fd_sc_hd__mux2_1 _3257_ (.A0(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[22] ),
    .A1(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[30] ),
    .S(_1222_),
    .X(_1366_));
 sky130_fd_sc_hd__a21oi_1 _3258_ (.A1(_1220_),
    .A2(_1366_),
    .B1(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_first_qq[2] ),
    .Y(_1367_));
 sky130_fd_sc_hd__a32o_1 _3259_ (.A1(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_first_qq[2] ),
    .A2(_1361_),
    .A3(_1363_),
    .B1(_1365_),
    .B2(_1367_),
    .X(_1368_));
 sky130_fd_sc_hd__a2bb2o_1 _3260_ (.A1_N(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_first_qq[3] ),
    .A2_N(_1368_),
    .B1(_1235_),
    .B2(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[70] ),
    .X(_1369_));
 sky130_fd_sc_hd__a32o_1 _3261_ (.A1(_1217_),
    .A2(_1334_),
    .A3(_1359_),
    .B1(_1369_),
    .B2(_0883_),
    .X(_1370_));
 sky130_fd_sc_hd__mux2_1 _3262_ (.A0(\usb2uart.u_usb_cdc.u_sie.rx_data[6] ),
    .A1(_1370_),
    .S(_1146_),
    .X(_1371_));
 sky130_fd_sc_hd__mux2_1 _3263_ (.A0(\usb2uart.u_usb_cdc.u_sie.data_q[6] ),
    .A1(_1371_),
    .S(_0836_),
    .X(_1372_));
 sky130_fd_sc_hd__clkbuf_1 _3264_ (.A(_1372_),
    .X(_0162_));
 sky130_fd_sc_hd__mux2_1 _3265_ (.A0(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[39] ),
    .A1(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[47] ),
    .S(_1223_),
    .X(_1373_));
 sky130_fd_sc_hd__or2b_1 _3266_ (.A(_1220_),
    .B_N(_1373_),
    .X(_1374_));
 sky130_fd_sc_hd__mux2_1 _3267_ (.A0(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[55] ),
    .A1(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[63] ),
    .S(_1261_),
    .X(_1375_));
 sky130_fd_sc_hd__nand2_1 _3268_ (.A(_1269_),
    .B(_1375_),
    .Y(_1376_));
 sky130_fd_sc_hd__mux2_1 _3269_ (.A0(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[7] ),
    .A1(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[15] ),
    .S(_1223_),
    .X(_1377_));
 sky130_fd_sc_hd__or2b_1 _3270_ (.A(_1221_),
    .B_N(_1377_),
    .X(_1378_));
 sky130_fd_sc_hd__mux2_1 _3271_ (.A0(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[23] ),
    .A1(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[31] ),
    .S(_1261_),
    .X(_1379_));
 sky130_fd_sc_hd__a21oi_1 _3272_ (.A1(_1269_),
    .A2(_1379_),
    .B1(_1227_),
    .Y(_1380_));
 sky130_fd_sc_hd__a32o_1 _3273_ (.A1(_1265_),
    .A2(_1374_),
    .A3(_1376_),
    .B1(_1378_),
    .B2(_1380_),
    .X(_1381_));
 sky130_fd_sc_hd__a2bb2o_1 _3274_ (.A1_N(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_first_qq[3] ),
    .A2_N(_1381_),
    .B1(_1235_),
    .B2(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[71] ),
    .X(_1382_));
 sky130_fd_sc_hd__a21oi_1 _3275_ (.A1(_1281_),
    .A2(_1342_),
    .B1(_1189_),
    .Y(_1383_));
 sky130_fd_sc_hd__a2111oi_1 _3276_ (.A1(_1240_),
    .A2(_2024_),
    .B1(\usb2uart.u_usb_cdc.u_ctrl_endp.byte_cnt_q[6] ),
    .C1(_1249_),
    .D1(_1383_),
    .Y(_1384_));
 sky130_fd_sc_hd__a221o_1 _3277_ (.A1(_0883_),
    .A2(_1382_),
    .B1(_1384_),
    .B2(_1216_),
    .C1(_0884_),
    .X(_1385_));
 sky130_fd_sc_hd__o21a_1 _3278_ (.A1(\usb2uart.u_usb_cdc.u_sie.rx_data[7] ),
    .A2(_1146_),
    .B1(_0836_),
    .X(_1386_));
 sky130_fd_sc_hd__a22o_1 _3279_ (.A1(\usb2uart.u_usb_cdc.u_sie.data_q[7] ),
    .A2(_0839_),
    .B1(_1385_),
    .B2(_1386_),
    .X(_0163_));
 sky130_fd_sc_hd__o21a_2 _3280_ (.A1(\usb2uart.u_usb_cdc.u_sie.phy_state_q[3] ),
    .A2(_0841_),
    .B1(_0591_),
    .X(_1387_));
 sky130_fd_sc_hd__a22o_1 _3281_ (.A1(_1119_),
    .A2(_0839_),
    .B1(_1387_),
    .B2(_0517_),
    .X(_0164_));
 sky130_fd_sc_hd__a22o_1 _3282_ (.A1(_1124_),
    .A2(_0839_),
    .B1(_1387_),
    .B2(_0521_),
    .X(_0165_));
 sky130_fd_sc_hd__a22o_1 _3283_ (.A1(_1126_),
    .A2(_0839_),
    .B1(_1387_),
    .B2(\usb2uart.u_usb_cdc.u_sie.data_q[2] ),
    .X(_0166_));
 sky130_fd_sc_hd__a22o_1 _3284_ (.A1(_1128_),
    .A2(_0839_),
    .B1(_1387_),
    .B2(_0519_),
    .X(_0167_));
 sky130_fd_sc_hd__a22o_1 _3285_ (.A1(_1130_),
    .A2(_0839_),
    .B1(_1387_),
    .B2(\usb2uart.u_usb_cdc.u_sie.data_q[4] ),
    .X(_0168_));
 sky130_fd_sc_hd__a22o_1 _3286_ (.A1(_1132_),
    .A2(_0839_),
    .B1(_1387_),
    .B2(\usb2uart.u_usb_cdc.u_sie.data_q[5] ),
    .X(_0169_));
 sky130_fd_sc_hd__a22o_1 _3287_ (.A1(_1134_),
    .A2(_0839_),
    .B1(_1387_),
    .B2(\usb2uart.u_usb_cdc.u_sie.data_q[6] ),
    .X(_0170_));
 sky130_fd_sc_hd__a22o_1 _3288_ (.A1(_1171_),
    .A2(_0839_),
    .B1(_1387_),
    .B2(\usb2uart.u_usb_cdc.u_sie.data_q[7] ),
    .X(_0171_));
 sky130_fd_sc_hd__a21o_2 _3289_ (.A1(_0688_),
    .A2(_0856_),
    .B1(_0690_),
    .X(_1388_));
 sky130_fd_sc_hd__mux2_1 _3290_ (.A0(_1119_),
    .A1(\usb2uart.u_usb_cdc.u_ctrl_endp.rec_q[0] ),
    .S(_1388_),
    .X(_1389_));
 sky130_fd_sc_hd__clkbuf_1 _3291_ (.A(_1389_),
    .X(_0172_));
 sky130_fd_sc_hd__mux2_1 _3292_ (.A0(_1124_),
    .A1(\usb2uart.u_usb_cdc.u_ctrl_endp.rec_q[1] ),
    .S(_1388_),
    .X(_1390_));
 sky130_fd_sc_hd__clkbuf_1 _3293_ (.A(_1390_),
    .X(_0173_));
 sky130_fd_sc_hd__or3_1 _3294_ (.A(_2081_),
    .B(_0488_),
    .C(_0498_),
    .X(_1391_));
 sky130_fd_sc_hd__a21o_1 _3295_ (.A1(_0473_),
    .A2(_0773_),
    .B1(_1391_),
    .X(_1392_));
 sky130_fd_sc_hd__mux2_1 _3296_ (.A0(_1171_),
    .A1(\usb2uart.u_usb_cdc.u_ctrl_endp.in_endp_q ),
    .S(_1392_),
    .X(_1393_));
 sky130_fd_sc_hd__clkbuf_1 _3297_ (.A(_1393_),
    .X(_0174_));
 sky130_fd_sc_hd__a31o_1 _3298_ (.A1(\usb2uart.u_usb_cdc.u_ctrl_endp.req_q[7] ),
    .A2(_0681_),
    .A3(_0858_),
    .B1(_0487_),
    .X(_1394_));
 sky130_fd_sc_hd__o21ba_1 _3299_ (.A1(_2012_),
    .A2(_1394_),
    .B1_N(_0690_),
    .X(_1395_));
 sky130_fd_sc_hd__mux2_1 _3300_ (.A0(\usb2uart.u_usb_cdc.u_ctrl_endp.dev_state_q[0] ),
    .A1(_0699_),
    .S(_1395_),
    .X(_1396_));
 sky130_fd_sc_hd__clkbuf_1 _3301_ (.A(_1396_),
    .X(_0175_));
 sky130_fd_sc_hd__or2_1 _3302_ (.A(\usb2uart.u_usb_cdc.u_ctrl_endp.dev_state_q[1] ),
    .B(_1395_),
    .X(_1397_));
 sky130_fd_sc_hd__clkbuf_1 _3303_ (.A(_1397_),
    .X(_0176_));
 sky130_fd_sc_hd__nor2_1 _3304_ (.A(_2075_),
    .B(_2005_),
    .Y(_1398_));
 sky130_fd_sc_hd__or2_1 _3305_ (.A(_0862_),
    .B(_1398_),
    .X(_1399_));
 sky130_fd_sc_hd__a22o_1 _3306_ (.A1(_0863_),
    .A2(_0865_),
    .B1(_1399_),
    .B2(\usb2uart.u_usb_cdc.bulk_out_nak ),
    .X(_0177_));
 sky130_fd_sc_hd__o31a_1 _3307_ (.A1(\usb2uart.u_usb_cdc.out_data[7] ),
    .A2(_0735_),
    .A3(_0489_),
    .B1(_0688_),
    .X(_1400_));
 sky130_fd_sc_hd__nor2_4 _3308_ (.A(_0690_),
    .B(_1400_),
    .Y(_1401_));
 sky130_fd_sc_hd__mux2_1 _3309_ (.A0(\usb2uart.u_usb_cdc.u_ctrl_endp.addr_q[0] ),
    .A1(_1119_),
    .S(_1401_),
    .X(_1402_));
 sky130_fd_sc_hd__clkbuf_1 _3310_ (.A(_1402_),
    .X(_0178_));
 sky130_fd_sc_hd__mux2_1 _3311_ (.A0(\usb2uart.u_usb_cdc.u_ctrl_endp.addr_q[1] ),
    .A1(_1124_),
    .S(_1401_),
    .X(_1403_));
 sky130_fd_sc_hd__clkbuf_1 _3312_ (.A(_1403_),
    .X(_0179_));
 sky130_fd_sc_hd__mux2_1 _3313_ (.A0(\usb2uart.u_usb_cdc.u_ctrl_endp.addr_q[2] ),
    .A1(_1126_),
    .S(_1401_),
    .X(_1404_));
 sky130_fd_sc_hd__clkbuf_1 _3314_ (.A(_1404_),
    .X(_0180_));
 sky130_fd_sc_hd__mux2_1 _3315_ (.A0(\usb2uart.u_usb_cdc.u_ctrl_endp.addr_q[3] ),
    .A1(_1128_),
    .S(_1401_),
    .X(_1405_));
 sky130_fd_sc_hd__clkbuf_1 _3316_ (.A(_1405_),
    .X(_0181_));
 sky130_fd_sc_hd__mux2_1 _3317_ (.A0(\usb2uart.u_usb_cdc.u_ctrl_endp.addr_q[4] ),
    .A1(_1130_),
    .S(_1401_),
    .X(_1406_));
 sky130_fd_sc_hd__clkbuf_1 _3318_ (.A(_1406_),
    .X(_0182_));
 sky130_fd_sc_hd__mux2_1 _3319_ (.A0(\usb2uart.u_usb_cdc.u_ctrl_endp.addr_q[5] ),
    .A1(_1132_),
    .S(_1401_),
    .X(_1407_));
 sky130_fd_sc_hd__clkbuf_1 _3320_ (.A(_1407_),
    .X(_0183_));
 sky130_fd_sc_hd__mux2_1 _3321_ (.A0(\usb2uart.u_usb_cdc.u_ctrl_endp.addr_q[6] ),
    .A1(_1134_),
    .S(_1401_),
    .X(_1408_));
 sky130_fd_sc_hd__clkbuf_1 _3322_ (.A(_1408_),
    .X(_0184_));
 sky130_fd_sc_hd__o31ai_1 _3323_ (.A1(_0645_),
    .A2(_2006_),
    .A3(_0655_),
    .B1(\usb2uart.u_usb_cdc.u_ctrl_endp.state_q[3] ),
    .Y(_1409_));
 sky130_fd_sc_hd__a21o_1 _3324_ (.A1(_2018_),
    .A2(_1409_),
    .B1(_2081_),
    .X(_1410_));
 sky130_fd_sc_hd__and3_2 _3325_ (.A(_2009_),
    .B(_2078_),
    .C(_1410_),
    .X(_1411_));
 sky130_fd_sc_hd__inv_2 _3326_ (.A(_1411_),
    .Y(_1412_));
 sky130_fd_sc_hd__o21ai_1 _3327_ (.A1(\usb2uart.u_usb_cdc.u_ctrl_endp.state_q[3] ),
    .A2(_0688_),
    .B1(_2020_),
    .Y(_1413_));
 sky130_fd_sc_hd__nor2_1 _3328_ (.A(_1412_),
    .B(_1413_),
    .Y(_1414_));
 sky130_fd_sc_hd__mux2_1 _3329_ (.A0(_1412_),
    .A1(_1414_),
    .S(_2084_),
    .X(_1415_));
 sky130_fd_sc_hd__clkbuf_1 _3330_ (.A(_1415_),
    .X(_0185_));
 sky130_fd_sc_hd__a32o_1 _3331_ (.A1(_0641_),
    .A2(_1242_),
    .A3(_1414_),
    .B1(_1412_),
    .B2(_0450_),
    .X(_0186_));
 sky130_fd_sc_hd__nor2_1 _3332_ (.A(_0502_),
    .B(_1241_),
    .Y(_1416_));
 sky130_fd_sc_hd__a22o_1 _3333_ (.A1(_1205_),
    .A2(_1412_),
    .B1(_1414_),
    .B2(_1416_),
    .X(_0187_));
 sky130_fd_sc_hd__nand3_1 _3334_ (.A(_1240_),
    .B(_0502_),
    .C(_1411_),
    .Y(_1417_));
 sky130_fd_sc_hd__nand2_1 _3335_ (.A(_1411_),
    .B(_1413_),
    .Y(_1418_));
 sky130_fd_sc_hd__a21o_1 _3336_ (.A1(_0502_),
    .A2(_1411_),
    .B1(_1240_),
    .X(_1419_));
 sky130_fd_sc_hd__and3_1 _3337_ (.A(_1417_),
    .B(_1418_),
    .C(_1419_),
    .X(_1420_));
 sky130_fd_sc_hd__clkbuf_1 _3338_ (.A(_1420_),
    .X(_0188_));
 sky130_fd_sc_hd__and4_1 _3339_ (.A(_1240_),
    .B(_1189_),
    .C(_0502_),
    .D(_1411_),
    .X(_1421_));
 sky130_fd_sc_hd__clkinv_2 _3340_ (.A(_1421_),
    .Y(_1422_));
 sky130_fd_sc_hd__a31o_1 _3341_ (.A1(_1240_),
    .A2(_0502_),
    .A3(_1411_),
    .B1(_1189_),
    .X(_1423_));
 sky130_fd_sc_hd__and3_1 _3342_ (.A(_1418_),
    .B(_1422_),
    .C(_1423_),
    .X(_1424_));
 sky130_fd_sc_hd__clkbuf_1 _3343_ (.A(_1424_),
    .X(_0189_));
 sky130_fd_sc_hd__and2_1 _3344_ (.A(_0454_),
    .B(_1421_),
    .X(_1425_));
 sky130_fd_sc_hd__o21ai_1 _3345_ (.A1(_0454_),
    .A2(_1421_),
    .B1(_1418_),
    .Y(_1426_));
 sky130_fd_sc_hd__nor2_1 _3346_ (.A(_1425_),
    .B(_1426_),
    .Y(_0190_));
 sky130_fd_sc_hd__a21boi_1 _3347_ (.A1(\usb2uart.u_usb_cdc.u_ctrl_endp.byte_cnt_q[6] ),
    .A2(_1425_),
    .B1_N(_1418_),
    .Y(_1427_));
 sky130_fd_sc_hd__o21a_1 _3348_ (.A1(\usb2uart.u_usb_cdc.u_ctrl_endp.byte_cnt_q[6] ),
    .A2(_1425_),
    .B1(_1427_),
    .X(_0191_));
 sky130_fd_sc_hd__o32a_1 _3349_ (.A1(_0485_),
    .A2(_0503_),
    .A3(_1309_),
    .B1(_0476_),
    .B2(_0506_),
    .X(_1428_));
 sky130_fd_sc_hd__a21oi_4 _3350_ (.A1(_0688_),
    .A2(_1428_),
    .B1(_0690_),
    .Y(_1429_));
 sky130_fd_sc_hd__o211ai_4 _3351_ (.A1(_0678_),
    .A2(_1309_),
    .B1(_1429_),
    .C1(_0503_),
    .Y(_1430_));
 sky130_fd_sc_hd__o22a_1 _3352_ (.A1(\usb2uart.u_usb_cdc.u_ctrl_endp.max_length_q[0] ),
    .A2(_1429_),
    .B1(_1430_),
    .B2(_1119_),
    .X(_0192_));
 sky130_fd_sc_hd__o22a_1 _3353_ (.A1(\usb2uart.u_usb_cdc.u_ctrl_endp.max_length_q[1] ),
    .A2(_1429_),
    .B1(_1430_),
    .B2(_1124_),
    .X(_0193_));
 sky130_fd_sc_hd__o22a_1 _3354_ (.A1(\usb2uart.u_usb_cdc.u_ctrl_endp.max_length_q[2] ),
    .A2(_1429_),
    .B1(_1430_),
    .B2(_1126_),
    .X(_0194_));
 sky130_fd_sc_hd__o22a_1 _3355_ (.A1(\usb2uart.u_usb_cdc.u_ctrl_endp.max_length_q[3] ),
    .A2(_1429_),
    .B1(_1430_),
    .B2(_1128_),
    .X(_0195_));
 sky130_fd_sc_hd__o22a_1 _3356_ (.A1(\usb2uart.u_usb_cdc.u_ctrl_endp.max_length_q[4] ),
    .A2(_1429_),
    .B1(_1430_),
    .B2(_1130_),
    .X(_0196_));
 sky130_fd_sc_hd__o22a_1 _3357_ (.A1(\usb2uart.u_usb_cdc.u_ctrl_endp.max_length_q[5] ),
    .A2(_1429_),
    .B1(_1430_),
    .B2(_1132_),
    .X(_0197_));
 sky130_fd_sc_hd__o22a_1 _3358_ (.A1(\usb2uart.u_usb_cdc.u_ctrl_endp.max_length_q[6] ),
    .A2(_1429_),
    .B1(_1430_),
    .B2(_1134_),
    .X(_0198_));
 sky130_fd_sc_hd__mux2_1 _3359_ (.A0(_1171_),
    .A1(_0461_),
    .S(_1388_),
    .X(_1431_));
 sky130_fd_sc_hd__clkbuf_1 _3360_ (.A(_1431_),
    .X(_0199_));
 sky130_fd_sc_hd__mux2_1 _3361_ (.A0(_1132_),
    .A1(\usb2uart.u_usb_cdc.u_ctrl_endp.class_q ),
    .S(_1388_),
    .X(_1432_));
 sky130_fd_sc_hd__clkbuf_1 _3362_ (.A(_1432_),
    .X(_0200_));
 sky130_fd_sc_hd__o31a_1 _3363_ (.A1(_0735_),
    .A2(_2017_),
    .A3(_0646_),
    .B1(_0473_),
    .X(_1433_));
 sky130_fd_sc_hd__nor2_4 _3364_ (.A(_1391_),
    .B(_1433_),
    .Y(_1434_));
 sky130_fd_sc_hd__mux2_1 _3365_ (.A0(\usb2uart.u_usb_cdc.addr[0] ),
    .A1(\usb2uart.u_usb_cdc.u_ctrl_endp.addr_q[0] ),
    .S(_1434_),
    .X(_1435_));
 sky130_fd_sc_hd__clkbuf_1 _3366_ (.A(_1435_),
    .X(_0201_));
 sky130_fd_sc_hd__mux2_1 _3367_ (.A0(\usb2uart.u_usb_cdc.addr[1] ),
    .A1(\usb2uart.u_usb_cdc.u_ctrl_endp.addr_q[1] ),
    .S(_1434_),
    .X(_1436_));
 sky130_fd_sc_hd__clkbuf_1 _3368_ (.A(_1436_),
    .X(_0202_));
 sky130_fd_sc_hd__mux2_1 _3369_ (.A0(\usb2uart.u_usb_cdc.addr[2] ),
    .A1(\usb2uart.u_usb_cdc.u_ctrl_endp.addr_q[2] ),
    .S(_1434_),
    .X(_1437_));
 sky130_fd_sc_hd__clkbuf_1 _3370_ (.A(_1437_),
    .X(_0203_));
 sky130_fd_sc_hd__mux2_1 _3371_ (.A0(\usb2uart.u_usb_cdc.addr[3] ),
    .A1(\usb2uart.u_usb_cdc.u_ctrl_endp.addr_q[3] ),
    .S(_1434_),
    .X(_1438_));
 sky130_fd_sc_hd__clkbuf_1 _3372_ (.A(_1438_),
    .X(_0204_));
 sky130_fd_sc_hd__mux2_1 _3373_ (.A0(\usb2uart.u_usb_cdc.addr[4] ),
    .A1(\usb2uart.u_usb_cdc.u_ctrl_endp.addr_q[4] ),
    .S(_1434_),
    .X(_1439_));
 sky130_fd_sc_hd__clkbuf_1 _3374_ (.A(_1439_),
    .X(_0205_));
 sky130_fd_sc_hd__mux2_1 _3375_ (.A0(\usb2uart.u_usb_cdc.addr[5] ),
    .A1(\usb2uart.u_usb_cdc.u_ctrl_endp.addr_q[5] ),
    .S(_1434_),
    .X(_1440_));
 sky130_fd_sc_hd__clkbuf_1 _3376_ (.A(_1440_),
    .X(_0206_));
 sky130_fd_sc_hd__mux2_1 _3377_ (.A0(\usb2uart.u_usb_cdc.addr[6] ),
    .A1(\usb2uart.u_usb_cdc.u_ctrl_endp.addr_q[6] ),
    .S(_1434_),
    .X(_1441_));
 sky130_fd_sc_hd__clkbuf_1 _3378_ (.A(_1441_),
    .X(_0207_));
 sky130_fd_sc_hd__buf_2 _3379_ (.A(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_last_qq[0] ),
    .X(_1442_));
 sky130_fd_sc_hd__buf_2 _3380_ (.A(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_last_qq[3] ),
    .X(_1443_));
 sky130_fd_sc_hd__or2_1 _3381_ (.A(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_last_qq[0] ),
    .B(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_last_qq[1] ),
    .X(_1444_));
 sky130_fd_sc_hd__nor2_1 _3382_ (.A(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_last_qq[2] ),
    .B(_1444_),
    .Y(_1445_));
 sky130_fd_sc_hd__nand2_1 _3383_ (.A(_1443_),
    .B(_1445_),
    .Y(_1446_));
 sky130_fd_sc_hd__nand2_1 _3384_ (.A(_2006_),
    .B(_1446_),
    .Y(_1447_));
 sky130_fd_sc_hd__mux2_1 _3385_ (.A0(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_last_qq[0] ),
    .A1(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_last_q[0] ),
    .S(\usb2uart.u_usb_cdc.bulk_out_nak ),
    .X(_1448_));
 sky130_fd_sc_hd__a2bb2o_1 _3386_ (.A1_N(_1442_),
    .A2_N(_1447_),
    .B1(_1448_),
    .B2(_0487_),
    .X(_1449_));
 sky130_fd_sc_hd__mux2_1 _3387_ (.A0(_1449_),
    .A1(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_last_q[0] ),
    .S(_0652_),
    .X(_1450_));
 sky130_fd_sc_hd__mux2_1 _3388_ (.A0(_1442_),
    .A1(_1450_),
    .S(_0866_),
    .X(_1451_));
 sky130_fd_sc_hd__clkbuf_1 _3389_ (.A(_1451_),
    .X(_0208_));
 sky130_fd_sc_hd__clkbuf_4 _3390_ (.A(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_last_qq[1] ),
    .X(_1452_));
 sky130_fd_sc_hd__mux2_1 _3391_ (.A0(_1452_),
    .A1(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_last_q[1] ),
    .S(\usb2uart.u_usb_cdc.bulk_out_nak ),
    .X(_1453_));
 sky130_fd_sc_hd__nand2_1 _3392_ (.A(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_last_qq[0] ),
    .B(_1452_),
    .Y(_1454_));
 sky130_fd_sc_hd__and3_1 _3393_ (.A(_2006_),
    .B(_1444_),
    .C(_1454_),
    .X(_1455_));
 sky130_fd_sc_hd__a21o_1 _3394_ (.A1(_0487_),
    .A2(_1453_),
    .B1(_1455_),
    .X(_1456_));
 sky130_fd_sc_hd__mux2_1 _3395_ (.A0(_1456_),
    .A1(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_last_q[1] ),
    .S(_0652_),
    .X(_1457_));
 sky130_fd_sc_hd__mux2_1 _3396_ (.A0(_1452_),
    .A1(_1457_),
    .S(_0866_),
    .X(_1458_));
 sky130_fd_sc_hd__clkbuf_1 _3397_ (.A(_1458_),
    .X(_0209_));
 sky130_fd_sc_hd__and3_2 _3398_ (.A(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_last_qq[0] ),
    .B(_1452_),
    .C(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_last_qq[2] ),
    .X(_1459_));
 sky130_fd_sc_hd__a21oi_1 _3399_ (.A1(_1442_),
    .A2(_1452_),
    .B1(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_last_qq[2] ),
    .Y(_1460_));
 sky130_fd_sc_hd__mux2_1 _3400_ (.A0(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_last_qq[2] ),
    .A1(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_last_q[2] ),
    .S(\usb2uart.u_usb_cdc.bulk_out_nak ),
    .X(_1461_));
 sky130_fd_sc_hd__a22oi_1 _3401_ (.A1(_0652_),
    .A2(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_last_q[2] ),
    .B1(_1398_),
    .B2(_1461_),
    .Y(_1462_));
 sky130_fd_sc_hd__o31a_1 _3402_ (.A1(_0661_),
    .A2(_1459_),
    .A3(_1460_),
    .B1(_1462_),
    .X(_1463_));
 sky130_fd_sc_hd__nand2_1 _3403_ (.A(_0866_),
    .B(_1463_),
    .Y(_1464_));
 sky130_fd_sc_hd__o21a_1 _3404_ (.A1(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_last_qq[2] ),
    .A2(_0866_),
    .B1(_1464_),
    .X(_0210_));
 sky130_fd_sc_hd__mux2_1 _3405_ (.A0(_1443_),
    .A1(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_last_q[3] ),
    .S(\usb2uart.u_usb_cdc.bulk_out_nak ),
    .X(_1465_));
 sky130_fd_sc_hd__o21bai_1 _3406_ (.A1(_1443_),
    .A2(_1459_),
    .B1_N(_2075_),
    .Y(_1466_));
 sky130_fd_sc_hd__a211oi_1 _3407_ (.A1(_1443_),
    .A2(_1459_),
    .B1(_1466_),
    .C1(_1447_),
    .Y(_1467_));
 sky130_fd_sc_hd__a221o_1 _3408_ (.A1(_0652_),
    .A2(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_last_q[3] ),
    .B1(_1398_),
    .B2(_1465_),
    .C1(_1467_),
    .X(_1468_));
 sky130_fd_sc_hd__mux2_1 _3409_ (.A0(_1443_),
    .A1(_1468_),
    .S(_0866_),
    .X(_1469_));
 sky130_fd_sc_hd__clkbuf_1 _3410_ (.A(_1469_),
    .X(_0211_));
 sky130_fd_sc_hd__nand2_2 _3411_ (.A(_0863_),
    .B(_1398_),
    .Y(_1470_));
 sky130_fd_sc_hd__mux2_1 _3412_ (.A0(_1448_),
    .A1(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_last_q[0] ),
    .S(_1470_),
    .X(_1471_));
 sky130_fd_sc_hd__clkbuf_1 _3413_ (.A(_1471_),
    .X(_0212_));
 sky130_fd_sc_hd__mux2_1 _3414_ (.A0(_1453_),
    .A1(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_last_q[1] ),
    .S(_1470_),
    .X(_1472_));
 sky130_fd_sc_hd__clkbuf_1 _3415_ (.A(_1472_),
    .X(_0213_));
 sky130_fd_sc_hd__mux2_1 _3416_ (.A0(_1461_),
    .A1(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_last_q[2] ),
    .S(_1470_),
    .X(_1473_));
 sky130_fd_sc_hd__clkbuf_1 _3417_ (.A(_1473_),
    .X(_0214_));
 sky130_fd_sc_hd__mux2_1 _3418_ (.A0(_1465_),
    .A1(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_last_q[3] ),
    .S(_1470_),
    .X(_1474_));
 sky130_fd_sc_hd__clkbuf_1 _3419_ (.A(_1474_),
    .X(_0215_));
 sky130_fd_sc_hd__or3_4 _3420_ (.A(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_last_qq[1] ),
    .B(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_last_qq[2] ),
    .C(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_last_qq[3] ),
    .X(_1475_));
 sky130_fd_sc_hd__or3_1 _3421_ (.A(_2075_),
    .B(_0864_),
    .C(_1399_),
    .X(_1476_));
 sky130_fd_sc_hd__or3_1 _3422_ (.A(_1442_),
    .B(_1475_),
    .C(_1476_),
    .X(_1477_));
 sky130_fd_sc_hd__clkbuf_4 _3423_ (.A(_1477_),
    .X(_1478_));
 sky130_fd_sc_hd__mux2_1 _3424_ (.A0(_1119_),
    .A1(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[0] ),
    .S(_1478_),
    .X(_1479_));
 sky130_fd_sc_hd__clkbuf_1 _3425_ (.A(_1479_),
    .X(_0216_));
 sky130_fd_sc_hd__mux2_1 _3426_ (.A0(_1124_),
    .A1(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[1] ),
    .S(_1478_),
    .X(_1480_));
 sky130_fd_sc_hd__clkbuf_1 _3427_ (.A(_1480_),
    .X(_0217_));
 sky130_fd_sc_hd__mux2_1 _3428_ (.A0(_1126_),
    .A1(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[2] ),
    .S(_1478_),
    .X(_1481_));
 sky130_fd_sc_hd__clkbuf_1 _3429_ (.A(_1481_),
    .X(_0218_));
 sky130_fd_sc_hd__mux2_1 _3430_ (.A0(_1128_),
    .A1(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[3] ),
    .S(_1478_),
    .X(_1482_));
 sky130_fd_sc_hd__clkbuf_1 _3431_ (.A(_1482_),
    .X(_0219_));
 sky130_fd_sc_hd__mux2_1 _3432_ (.A0(_1130_),
    .A1(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[4] ),
    .S(_1478_),
    .X(_1483_));
 sky130_fd_sc_hd__clkbuf_1 _3433_ (.A(_1483_),
    .X(_0220_));
 sky130_fd_sc_hd__mux2_1 _3434_ (.A0(_1132_),
    .A1(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[5] ),
    .S(_1478_),
    .X(_1484_));
 sky130_fd_sc_hd__clkbuf_1 _3435_ (.A(_1484_),
    .X(_0221_));
 sky130_fd_sc_hd__mux2_1 _3436_ (.A0(_1134_),
    .A1(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[6] ),
    .S(_1478_),
    .X(_1485_));
 sky130_fd_sc_hd__clkbuf_1 _3437_ (.A(_1485_),
    .X(_0222_));
 sky130_fd_sc_hd__mux2_1 _3438_ (.A0(_1171_),
    .A1(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[7] ),
    .S(_1478_),
    .X(_1486_));
 sky130_fd_sc_hd__clkbuf_1 _3439_ (.A(_1486_),
    .X(_0223_));
 sky130_fd_sc_hd__or3_1 _3440_ (.A(_2075_),
    .B(_0864_),
    .C(_1399_),
    .X(_1487_));
 sky130_fd_sc_hd__or3_1 _3441_ (.A(_1443_),
    .B(_1445_),
    .C(_1487_),
    .X(_1488_));
 sky130_fd_sc_hd__nor3_4 _3442_ (.A(_1452_),
    .B(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_last_qq[2] ),
    .C(_1488_),
    .Y(_1489_));
 sky130_fd_sc_hd__mux2_1 _3443_ (.A0(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[8] ),
    .A1(_1119_),
    .S(_1489_),
    .X(_1490_));
 sky130_fd_sc_hd__clkbuf_1 _3444_ (.A(_1490_),
    .X(_0224_));
 sky130_fd_sc_hd__mux2_1 _3445_ (.A0(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[9] ),
    .A1(_1124_),
    .S(_1489_),
    .X(_1491_));
 sky130_fd_sc_hd__clkbuf_1 _3446_ (.A(_1491_),
    .X(_0225_));
 sky130_fd_sc_hd__mux2_1 _3447_ (.A0(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[10] ),
    .A1(_1126_),
    .S(_1489_),
    .X(_1492_));
 sky130_fd_sc_hd__clkbuf_1 _3448_ (.A(_1492_),
    .X(_0226_));
 sky130_fd_sc_hd__mux2_1 _3449_ (.A0(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[11] ),
    .A1(_1128_),
    .S(_1489_),
    .X(_1493_));
 sky130_fd_sc_hd__clkbuf_1 _3450_ (.A(_1493_),
    .X(_0227_));
 sky130_fd_sc_hd__mux2_1 _3451_ (.A0(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[12] ),
    .A1(_1130_),
    .S(_1489_),
    .X(_1494_));
 sky130_fd_sc_hd__clkbuf_1 _3452_ (.A(_1494_),
    .X(_0228_));
 sky130_fd_sc_hd__mux2_1 _3453_ (.A0(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[13] ),
    .A1(_1132_),
    .S(_1489_),
    .X(_1495_));
 sky130_fd_sc_hd__clkbuf_1 _3454_ (.A(_1495_),
    .X(_0229_));
 sky130_fd_sc_hd__mux2_1 _3455_ (.A0(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[14] ),
    .A1(_1134_),
    .S(_1489_),
    .X(_1496_));
 sky130_fd_sc_hd__clkbuf_1 _3456_ (.A(_1496_),
    .X(_0230_));
 sky130_fd_sc_hd__mux2_1 _3457_ (.A0(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[15] ),
    .A1(_1171_),
    .S(_1489_),
    .X(_1497_));
 sky130_fd_sc_hd__clkbuf_1 _3458_ (.A(_1497_),
    .X(_0231_));
 sky130_fd_sc_hd__and2_1 _3459_ (.A(_0482_),
    .B(_1475_),
    .X(_1498_));
 sky130_fd_sc_hd__or3_1 _3460_ (.A(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_last_qq[3] ),
    .B(_1445_),
    .C(_1476_),
    .X(_1499_));
 sky130_fd_sc_hd__nand2_1 _3461_ (.A(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_last_qq[2] ),
    .B(_1444_),
    .Y(_1500_));
 sky130_fd_sc_hd__or2b_2 _3462_ (.A(_1499_),
    .B_N(_1500_),
    .X(_1501_));
 sky130_fd_sc_hd__nor3b_4 _3463_ (.A(_1501_),
    .B(_1442_),
    .C_N(_1452_),
    .Y(_1502_));
 sky130_fd_sc_hd__mux2_1 _3464_ (.A0(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[16] ),
    .A1(_1498_),
    .S(_1502_),
    .X(_1503_));
 sky130_fd_sc_hd__clkbuf_1 _3465_ (.A(_1503_),
    .X(_0232_));
 sky130_fd_sc_hd__and2_1 _3466_ (.A(_0465_),
    .B(_1475_),
    .X(_1504_));
 sky130_fd_sc_hd__mux2_1 _3467_ (.A0(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[17] ),
    .A1(_1504_),
    .S(_1502_),
    .X(_1505_));
 sky130_fd_sc_hd__clkbuf_1 _3468_ (.A(_1505_),
    .X(_0233_));
 sky130_fd_sc_hd__and2_1 _3469_ (.A(\usb2uart.u_usb_cdc.out_data[2] ),
    .B(_1475_),
    .X(_1506_));
 sky130_fd_sc_hd__mux2_1 _3470_ (.A0(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[18] ),
    .A1(_1506_),
    .S(_1502_),
    .X(_1507_));
 sky130_fd_sc_hd__clkbuf_1 _3471_ (.A(_1507_),
    .X(_0234_));
 sky130_fd_sc_hd__and2_1 _3472_ (.A(\usb2uart.u_usb_cdc.out_data[3] ),
    .B(_1475_),
    .X(_1508_));
 sky130_fd_sc_hd__mux2_1 _3473_ (.A0(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[19] ),
    .A1(_1508_),
    .S(_1502_),
    .X(_1509_));
 sky130_fd_sc_hd__clkbuf_1 _3474_ (.A(_1509_),
    .X(_0235_));
 sky130_fd_sc_hd__and2_1 _3475_ (.A(\usb2uart.u_usb_cdc.out_data[4] ),
    .B(_1475_),
    .X(_1510_));
 sky130_fd_sc_hd__mux2_1 _3476_ (.A0(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[20] ),
    .A1(_1510_),
    .S(_1502_),
    .X(_1511_));
 sky130_fd_sc_hd__clkbuf_1 _3477_ (.A(_1511_),
    .X(_0236_));
 sky130_fd_sc_hd__and2_1 _3478_ (.A(\usb2uart.u_usb_cdc.out_data[5] ),
    .B(_1475_),
    .X(_1512_));
 sky130_fd_sc_hd__mux2_1 _3479_ (.A0(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[21] ),
    .A1(_1512_),
    .S(_1502_),
    .X(_1513_));
 sky130_fd_sc_hd__clkbuf_1 _3480_ (.A(_1513_),
    .X(_0237_));
 sky130_fd_sc_hd__mux2_1 _3481_ (.A0(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[22] ),
    .A1(_1134_),
    .S(_1502_),
    .X(_1514_));
 sky130_fd_sc_hd__clkbuf_1 _3482_ (.A(_1514_),
    .X(_0238_));
 sky130_fd_sc_hd__mux2_1 _3483_ (.A0(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[23] ),
    .A1(_1171_),
    .S(_1502_),
    .X(_1515_));
 sky130_fd_sc_hd__clkbuf_1 _3484_ (.A(_1515_),
    .X(_0239_));
 sky130_fd_sc_hd__nor2_4 _3485_ (.A(_1454_),
    .B(_1501_),
    .Y(_1516_));
 sky130_fd_sc_hd__mux2_1 _3486_ (.A0(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[24] ),
    .A1(_1119_),
    .S(_1516_),
    .X(_1517_));
 sky130_fd_sc_hd__clkbuf_1 _3487_ (.A(_1517_),
    .X(_0240_));
 sky130_fd_sc_hd__mux2_1 _3488_ (.A0(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[25] ),
    .A1(_1124_),
    .S(_1516_),
    .X(_1518_));
 sky130_fd_sc_hd__clkbuf_1 _3489_ (.A(_1518_),
    .X(_0241_));
 sky130_fd_sc_hd__mux2_1 _3490_ (.A0(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[26] ),
    .A1(_1126_),
    .S(_1516_),
    .X(_1519_));
 sky130_fd_sc_hd__clkbuf_1 _3491_ (.A(_1519_),
    .X(_0242_));
 sky130_fd_sc_hd__mux2_1 _3492_ (.A0(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[27] ),
    .A1(_1128_),
    .S(_1516_),
    .X(_1520_));
 sky130_fd_sc_hd__clkbuf_1 _3493_ (.A(_1520_),
    .X(_0243_));
 sky130_fd_sc_hd__mux2_1 _3494_ (.A0(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[28] ),
    .A1(_1130_),
    .S(_1516_),
    .X(_1521_));
 sky130_fd_sc_hd__clkbuf_1 _3495_ (.A(_1521_),
    .X(_0244_));
 sky130_fd_sc_hd__mux2_1 _3496_ (.A0(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[29] ),
    .A1(_1132_),
    .S(_1516_),
    .X(_1522_));
 sky130_fd_sc_hd__clkbuf_1 _3497_ (.A(_1522_),
    .X(_0245_));
 sky130_fd_sc_hd__mux2_1 _3498_ (.A0(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[30] ),
    .A1(_0466_),
    .S(_1516_),
    .X(_1523_));
 sky130_fd_sc_hd__clkbuf_1 _3499_ (.A(_1523_),
    .X(_0246_));
 sky130_fd_sc_hd__mux2_1 _3500_ (.A0(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[31] ),
    .A1(\usb2uart.u_usb_cdc.out_data[7] ),
    .S(_1516_),
    .X(_1524_));
 sky130_fd_sc_hd__clkbuf_1 _3501_ (.A(_1524_),
    .X(_0247_));
 sky130_fd_sc_hd__or2_1 _3502_ (.A(_1444_),
    .B(_1499_),
    .X(_1525_));
 sky130_fd_sc_hd__buf_4 _3503_ (.A(_1525_),
    .X(_1526_));
 sky130_fd_sc_hd__mux2_1 _3504_ (.A0(_1498_),
    .A1(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[32] ),
    .S(_1526_),
    .X(_1527_));
 sky130_fd_sc_hd__clkbuf_1 _3505_ (.A(_1527_),
    .X(_0248_));
 sky130_fd_sc_hd__mux2_1 _3506_ (.A0(_1504_),
    .A1(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[33] ),
    .S(_1526_),
    .X(_1528_));
 sky130_fd_sc_hd__clkbuf_1 _3507_ (.A(_1528_),
    .X(_0249_));
 sky130_fd_sc_hd__mux2_1 _3508_ (.A0(_1506_),
    .A1(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[34] ),
    .S(_1526_),
    .X(_1529_));
 sky130_fd_sc_hd__clkbuf_1 _3509_ (.A(_1529_),
    .X(_0250_));
 sky130_fd_sc_hd__mux2_1 _3510_ (.A0(_1508_),
    .A1(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[35] ),
    .S(_1526_),
    .X(_1530_));
 sky130_fd_sc_hd__clkbuf_1 _3511_ (.A(_1530_),
    .X(_0251_));
 sky130_fd_sc_hd__mux2_1 _3512_ (.A0(_1510_),
    .A1(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[36] ),
    .S(_1526_),
    .X(_1531_));
 sky130_fd_sc_hd__clkbuf_1 _3513_ (.A(_1531_),
    .X(_0252_));
 sky130_fd_sc_hd__mux2_1 _3514_ (.A0(_1512_),
    .A1(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[37] ),
    .S(_1526_),
    .X(_1532_));
 sky130_fd_sc_hd__clkbuf_1 _3515_ (.A(_1532_),
    .X(_0253_));
 sky130_fd_sc_hd__mux2_1 _3516_ (.A0(_1134_),
    .A1(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[38] ),
    .S(_1526_),
    .X(_1533_));
 sky130_fd_sc_hd__clkbuf_1 _3517_ (.A(_1533_),
    .X(_0254_));
 sky130_fd_sc_hd__mux2_1 _3518_ (.A0(_1171_),
    .A1(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[39] ),
    .S(_1526_),
    .X(_1534_));
 sky130_fd_sc_hd__clkbuf_1 _3519_ (.A(_1534_),
    .X(_0255_));
 sky130_fd_sc_hd__or2_1 _3520_ (.A(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_last_qq[3] ),
    .B(_1500_),
    .X(_1535_));
 sky130_fd_sc_hd__or4b_1 _3521_ (.A(_1452_),
    .B(_1476_),
    .C(_1535_),
    .D_N(_1442_),
    .X(_1536_));
 sky130_fd_sc_hd__clkbuf_4 _3522_ (.A(_1536_),
    .X(_1537_));
 sky130_fd_sc_hd__mux2_1 _3523_ (.A0(_1119_),
    .A1(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[40] ),
    .S(_1537_),
    .X(_1538_));
 sky130_fd_sc_hd__clkbuf_1 _3524_ (.A(_1538_),
    .X(_0256_));
 sky130_fd_sc_hd__mux2_1 _3525_ (.A0(_1124_),
    .A1(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[41] ),
    .S(_1537_),
    .X(_1539_));
 sky130_fd_sc_hd__clkbuf_1 _3526_ (.A(_1539_),
    .X(_0257_));
 sky130_fd_sc_hd__mux2_1 _3527_ (.A0(_1126_),
    .A1(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[42] ),
    .S(_1537_),
    .X(_1540_));
 sky130_fd_sc_hd__clkbuf_1 _3528_ (.A(_1540_),
    .X(_0258_));
 sky130_fd_sc_hd__mux2_1 _3529_ (.A0(_1128_),
    .A1(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[43] ),
    .S(_1537_),
    .X(_1541_));
 sky130_fd_sc_hd__clkbuf_1 _3530_ (.A(_1541_),
    .X(_0259_));
 sky130_fd_sc_hd__mux2_1 _3531_ (.A0(_1130_),
    .A1(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[44] ),
    .S(_1537_),
    .X(_1542_));
 sky130_fd_sc_hd__clkbuf_1 _3532_ (.A(_1542_),
    .X(_0260_));
 sky130_fd_sc_hd__mux2_1 _3533_ (.A0(_1132_),
    .A1(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[45] ),
    .S(_1537_),
    .X(_1543_));
 sky130_fd_sc_hd__clkbuf_1 _3534_ (.A(_1543_),
    .X(_0261_));
 sky130_fd_sc_hd__mux2_1 _3535_ (.A0(_1134_),
    .A1(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[46] ),
    .S(_1537_),
    .X(_1544_));
 sky130_fd_sc_hd__clkbuf_1 _3536_ (.A(_1544_),
    .X(_0262_));
 sky130_fd_sc_hd__mux2_1 _3537_ (.A0(_1171_),
    .A1(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[47] ),
    .S(_1537_),
    .X(_1545_));
 sky130_fd_sc_hd__clkbuf_1 _3538_ (.A(_1545_),
    .X(_0263_));
 sky130_fd_sc_hd__or3_2 _3539_ (.A(_0661_),
    .B(_0862_),
    .C(_0864_),
    .X(_1546_));
 sky130_fd_sc_hd__or4_1 _3540_ (.A(_1442_),
    .B(_1443_),
    .C(_1546_),
    .D(_1500_),
    .X(_1547_));
 sky130_fd_sc_hd__clkbuf_4 _3541_ (.A(_1547_),
    .X(_1548_));
 sky130_fd_sc_hd__mux2_1 _3542_ (.A0(_1498_),
    .A1(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[48] ),
    .S(_1548_),
    .X(_1549_));
 sky130_fd_sc_hd__clkbuf_1 _3543_ (.A(_1549_),
    .X(_0264_));
 sky130_fd_sc_hd__mux2_1 _3544_ (.A0(_1504_),
    .A1(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[49] ),
    .S(_1548_),
    .X(_1550_));
 sky130_fd_sc_hd__clkbuf_1 _3545_ (.A(_1550_),
    .X(_0265_));
 sky130_fd_sc_hd__mux2_1 _3546_ (.A0(_1506_),
    .A1(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[50] ),
    .S(_1548_),
    .X(_1551_));
 sky130_fd_sc_hd__clkbuf_1 _3547_ (.A(_1551_),
    .X(_0266_));
 sky130_fd_sc_hd__mux2_1 _3548_ (.A0(_1508_),
    .A1(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[51] ),
    .S(_1548_),
    .X(_1552_));
 sky130_fd_sc_hd__clkbuf_1 _3549_ (.A(_1552_),
    .X(_0267_));
 sky130_fd_sc_hd__mux2_1 _3550_ (.A0(_1510_),
    .A1(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[52] ),
    .S(_1548_),
    .X(_1553_));
 sky130_fd_sc_hd__clkbuf_1 _3551_ (.A(_1553_),
    .X(_0268_));
 sky130_fd_sc_hd__mux2_1 _3552_ (.A0(_1512_),
    .A1(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[53] ),
    .S(_1548_),
    .X(_1554_));
 sky130_fd_sc_hd__clkbuf_1 _3553_ (.A(_1554_),
    .X(_0269_));
 sky130_fd_sc_hd__and2_1 _3554_ (.A(_0466_),
    .B(_1475_),
    .X(_1555_));
 sky130_fd_sc_hd__mux2_1 _3555_ (.A0(_1555_),
    .A1(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[54] ),
    .S(_1548_),
    .X(_1556_));
 sky130_fd_sc_hd__clkbuf_1 _3556_ (.A(_1556_),
    .X(_0270_));
 sky130_fd_sc_hd__and2_1 _3557_ (.A(\usb2uart.u_usb_cdc.out_data[7] ),
    .B(_1475_),
    .X(_1557_));
 sky130_fd_sc_hd__mux2_1 _3558_ (.A0(_1557_),
    .A1(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[55] ),
    .S(_1548_),
    .X(_1558_));
 sky130_fd_sc_hd__clkbuf_1 _3559_ (.A(_1558_),
    .X(_0271_));
 sky130_fd_sc_hd__nor2_1 _3560_ (.A(_1443_),
    .B(_1546_),
    .Y(_1559_));
 sky130_fd_sc_hd__nand2_4 _3561_ (.A(_1459_),
    .B(_1559_),
    .Y(_1560_));
 sky130_fd_sc_hd__and3_1 _3562_ (.A(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_last_qq[2] ),
    .B(_1444_),
    .C(_1559_),
    .X(_1561_));
 sky130_fd_sc_hd__and3_1 _3563_ (.A(_1442_),
    .B(_1452_),
    .C(_1561_),
    .X(_1562_));
 sky130_fd_sc_hd__buf_2 _3564_ (.A(_1562_),
    .X(_1563_));
 sky130_fd_sc_hd__a22o_1 _3565_ (.A1(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[56] ),
    .A2(_1560_),
    .B1(_1563_),
    .B2(_1119_),
    .X(_0272_));
 sky130_fd_sc_hd__a22o_1 _3566_ (.A1(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[57] ),
    .A2(_1560_),
    .B1(_1563_),
    .B2(_1124_),
    .X(_0273_));
 sky130_fd_sc_hd__a22o_1 _3567_ (.A1(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[58] ),
    .A2(_1560_),
    .B1(_1563_),
    .B2(_1126_),
    .X(_0274_));
 sky130_fd_sc_hd__a22o_1 _3568_ (.A1(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[59] ),
    .A2(_1560_),
    .B1(_1563_),
    .B2(_1128_),
    .X(_0275_));
 sky130_fd_sc_hd__a22o_1 _3569_ (.A1(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[60] ),
    .A2(_1560_),
    .B1(_1563_),
    .B2(_1130_),
    .X(_0276_));
 sky130_fd_sc_hd__a22o_1 _3570_ (.A1(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[61] ),
    .A2(_1560_),
    .B1(_1563_),
    .B2(_1132_),
    .X(_0277_));
 sky130_fd_sc_hd__a22o_1 _3571_ (.A1(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[62] ),
    .A2(_1560_),
    .B1(_1563_),
    .B2(_1134_),
    .X(_0278_));
 sky130_fd_sc_hd__a22o_1 _3572_ (.A1(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[63] ),
    .A2(_1560_),
    .B1(_1563_),
    .B2(_1171_),
    .X(_0279_));
 sky130_fd_sc_hd__nor2_4 _3573_ (.A(_1446_),
    .B(_1546_),
    .Y(_1564_));
 sky130_fd_sc_hd__mux2_1 _3574_ (.A0(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[64] ),
    .A1(_0482_),
    .S(_1564_),
    .X(_1565_));
 sky130_fd_sc_hd__clkbuf_1 _3575_ (.A(_1565_),
    .X(_0280_));
 sky130_fd_sc_hd__mux2_1 _3576_ (.A0(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[65] ),
    .A1(_0465_),
    .S(_1564_),
    .X(_1566_));
 sky130_fd_sc_hd__clkbuf_1 _3577_ (.A(_1566_),
    .X(_0281_));
 sky130_fd_sc_hd__mux2_1 _3578_ (.A0(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[66] ),
    .A1(_1126_),
    .S(_1564_),
    .X(_1567_));
 sky130_fd_sc_hd__clkbuf_1 _3579_ (.A(_1567_),
    .X(_0282_));
 sky130_fd_sc_hd__mux2_1 _3580_ (.A0(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[67] ),
    .A1(_1128_),
    .S(_1564_),
    .X(_1568_));
 sky130_fd_sc_hd__clkbuf_1 _3581_ (.A(_1568_),
    .X(_0283_));
 sky130_fd_sc_hd__mux2_1 _3582_ (.A0(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[68] ),
    .A1(_1130_),
    .S(_1564_),
    .X(_1569_));
 sky130_fd_sc_hd__clkbuf_1 _3583_ (.A(_1569_),
    .X(_0284_));
 sky130_fd_sc_hd__mux2_1 _3584_ (.A0(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[69] ),
    .A1(\usb2uart.u_usb_cdc.out_data[5] ),
    .S(_1564_),
    .X(_1570_));
 sky130_fd_sc_hd__clkbuf_1 _3585_ (.A(_1570_),
    .X(_0285_));
 sky130_fd_sc_hd__mux2_1 _3586_ (.A0(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[70] ),
    .A1(_0466_),
    .S(_1564_),
    .X(_1571_));
 sky130_fd_sc_hd__clkbuf_1 _3587_ (.A(_1571_),
    .X(_0286_));
 sky130_fd_sc_hd__mux2_1 _3588_ (.A0(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[71] ),
    .A1(\usb2uart.u_usb_cdc.out_data[7] ),
    .S(_1564_),
    .X(_1572_));
 sky130_fd_sc_hd__clkbuf_1 _3589_ (.A(_1572_),
    .X(_0287_));
 sky130_fd_sc_hd__inv_2 _3590_ (.A(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.delay_out_cnt_q[1] ),
    .Y(_1573_));
 sky130_fd_sc_hd__xor2_1 _3591_ (.A(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_last_q[1] ),
    .B(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_first_q[1] ),
    .X(_1574_));
 sky130_fd_sc_hd__xor2_1 _3592_ (.A(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_last_q[0] ),
    .B(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_first_q[0] ),
    .X(_1575_));
 sky130_fd_sc_hd__xor2_1 _3593_ (.A(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_last_q[3] ),
    .B(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_first_q[3] ),
    .X(_1576_));
 sky130_fd_sc_hd__xor2_1 _3594_ (.A(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_last_q[2] ),
    .B(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_first_q[2] ),
    .X(_1577_));
 sky130_fd_sc_hd__or4_1 _3595_ (.A(_1574_),
    .B(_1575_),
    .C(_1576_),
    .D(_1577_),
    .X(_1578_));
 sky130_fd_sc_hd__and2_1 _3596_ (.A(\usb2uart.u_uart.uart_tx_inst.s_axis_tready_reg ),
    .B(_1578_),
    .X(_1579_));
 sky130_fd_sc_hd__o21ai_1 _3597_ (.A1(_1573_),
    .A2(_1579_),
    .B1(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.delay_out_cnt_q[0] ),
    .Y(_0288_));
 sky130_fd_sc_hd__and3_1 _3598_ (.A(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.delay_out_cnt_q[1] ),
    .B(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.delay_out_cnt_q[0] ),
    .C(_1579_),
    .X(_1580_));
 sky130_fd_sc_hd__o21ba_1 _3599_ (.A1(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.delay_out_cnt_q[1] ),
    .A2(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.delay_out_cnt_q[0] ),
    .B1_N(_1580_),
    .X(_0289_));
 sky130_fd_sc_hd__xor2_1 _3600_ (.A(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_last_q[1] ),
    .B(_1260_),
    .X(_1581_));
 sky130_fd_sc_hd__buf_2 _3601_ (.A(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_last_q[0] ),
    .X(_1582_));
 sky130_fd_sc_hd__xor2_1 _3602_ (.A(_1582_),
    .B(_1267_),
    .X(_1583_));
 sky130_fd_sc_hd__xor2_1 _3603_ (.A(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_last_q[2] ),
    .B(_1265_),
    .X(_1584_));
 sky130_fd_sc_hd__xor2_1 _3604_ (.A(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_last_q[3] ),
    .B(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_first_qq[3] ),
    .X(_1585_));
 sky130_fd_sc_hd__or4_1 _3605_ (.A(_1581_),
    .B(_1583_),
    .C(_1584_),
    .D(_1585_),
    .X(_1586_));
 sky130_fd_sc_hd__nor2_1 _3606_ (.A(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_req_q ),
    .B(_0779_),
    .Y(_1587_));
 sky130_fd_sc_hd__xor2_1 _3607_ (.A(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_first_q[3] ),
    .B(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_last_q[3] ),
    .X(_1588_));
 sky130_fd_sc_hd__buf_2 _3608_ (.A(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_last_q[1] ),
    .X(_1589_));
 sky130_fd_sc_hd__xor2_1 _3609_ (.A(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_first_q[1] ),
    .B(_1589_),
    .X(_1590_));
 sky130_fd_sc_hd__xor2_1 _3610_ (.A(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_last_q[0] ),
    .B(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_first_q[0] ),
    .X(_1591_));
 sky130_fd_sc_hd__xor2_1 _3611_ (.A(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_first_q[2] ),
    .B(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_last_q[2] ),
    .X(_1592_));
 sky130_fd_sc_hd__or4_1 _3612_ (.A(_1588_),
    .B(_1590_),
    .C(_1591_),
    .D(_1592_),
    .X(_1593_));
 sky130_fd_sc_hd__a32o_1 _3613_ (.A1(\usb2uart.u_usb_cdc.bulk_in_valid ),
    .A2(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_req_q ),
    .A3(_1586_),
    .B1(_1587_),
    .B2(_1593_),
    .X(_0290_));
 sky130_fd_sc_hd__buf_4 _3614_ (.A(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_first_q[0] ),
    .X(_1594_));
 sky130_fd_sc_hd__buf_2 _3615_ (.A(_1594_),
    .X(_1595_));
 sky130_fd_sc_hd__and2_1 _3616_ (.A(_1595_),
    .B(_1580_),
    .X(_1596_));
 sky130_fd_sc_hd__inv_2 _3617_ (.A(_1596_),
    .Y(_1597_));
 sky130_fd_sc_hd__buf_2 _3618_ (.A(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_first_q[1] ),
    .X(_1598_));
 sky130_fd_sc_hd__or2_1 _3619_ (.A(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_first_q[0] ),
    .B(_1598_),
    .X(_1599_));
 sky130_fd_sc_hd__inv_2 _3620_ (.A(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_first_q[2] ),
    .Y(_1600_));
 sky130_fd_sc_hd__and3b_1 _3621_ (.A_N(_1599_),
    .B(_1600_),
    .C(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_first_q[3] ),
    .X(_1601_));
 sky130_fd_sc_hd__clkbuf_4 _3622_ (.A(_1601_),
    .X(_1602_));
 sky130_fd_sc_hd__nand2_1 _3623_ (.A(_1580_),
    .B(_1602_),
    .Y(_1603_));
 sky130_fd_sc_hd__o211a_1 _3624_ (.A1(_1595_),
    .A2(_1580_),
    .B1(_1597_),
    .C1(_1603_),
    .X(_0291_));
 sky130_fd_sc_hd__buf_2 _3625_ (.A(_1598_),
    .X(_1604_));
 sky130_fd_sc_hd__buf_2 _3626_ (.A(_1604_),
    .X(_1605_));
 sky130_fd_sc_hd__nand2_1 _3627_ (.A(_1605_),
    .B(_1596_),
    .Y(_1606_));
 sky130_fd_sc_hd__or2_1 _3628_ (.A(_1605_),
    .B(_1596_),
    .X(_1607_));
 sky130_fd_sc_hd__and2_1 _3629_ (.A(_1606_),
    .B(_1607_),
    .X(_1608_));
 sky130_fd_sc_hd__clkbuf_1 _3630_ (.A(_1608_),
    .X(_0292_));
 sky130_fd_sc_hd__clkbuf_4 _3631_ (.A(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_first_q[2] ),
    .X(_1609_));
 sky130_fd_sc_hd__xnor2_1 _3632_ (.A(_1609_),
    .B(_1606_),
    .Y(_0293_));
 sky130_fd_sc_hd__clkbuf_4 _3633_ (.A(_1600_),
    .X(_1610_));
 sky130_fd_sc_hd__inv_2 _3634_ (.A(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_first_q[3] ),
    .Y(_1611_));
 sky130_fd_sc_hd__a31o_1 _3635_ (.A1(_1605_),
    .A2(_1609_),
    .A3(_1596_),
    .B1(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_first_q[3] ),
    .X(_1612_));
 sky130_fd_sc_hd__o311a_1 _3636_ (.A1(_1610_),
    .A2(_1611_),
    .A3(_1606_),
    .B1(_1612_),
    .C1(_1603_),
    .X(_0294_));
 sky130_fd_sc_hd__and3b_1 _3637_ (.A_N(_1599_),
    .B(_1611_),
    .C(_1610_),
    .X(_1613_));
 sky130_fd_sc_hd__or3_1 _3638_ (.A(_1595_),
    .B(_1442_),
    .C(_1613_),
    .X(_1614_));
 sky130_fd_sc_hd__nand2_1 _3639_ (.A(_1595_),
    .B(_1605_),
    .Y(_1615_));
 sky130_fd_sc_hd__a21oi_1 _3640_ (.A1(_1599_),
    .A2(_1615_),
    .B1(_1613_),
    .Y(_1616_));
 sky130_fd_sc_hd__xnor2_1 _3641_ (.A(_1452_),
    .B(_1616_),
    .Y(_1617_));
 sky130_fd_sc_hd__o21a_1 _3642_ (.A1(_1609_),
    .A2(_1599_),
    .B1(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_first_q[3] ),
    .X(_1618_));
 sky130_fd_sc_hd__o21ai_1 _3643_ (.A1(_1613_),
    .A2(_1618_),
    .B1(_1443_),
    .Y(_1619_));
 sky130_fd_sc_hd__or3_1 _3644_ (.A(_1443_),
    .B(_1613_),
    .C(_1618_),
    .X(_1620_));
 sky130_fd_sc_hd__a21oi_1 _3645_ (.A1(_1609_),
    .A2(_1599_),
    .B1(_1602_),
    .Y(_1621_));
 sky130_fd_sc_hd__xnor2_1 _3646_ (.A(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_last_qq[2] ),
    .B(_1621_),
    .Y(_1622_));
 sky130_fd_sc_hd__o21a_1 _3647_ (.A1(_1595_),
    .A2(_1613_),
    .B1(_1442_),
    .X(_1623_));
 sky130_fd_sc_hd__nand2_1 _3648_ (.A(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.delay_out_cnt_q[1] ),
    .B(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.delay_out_cnt_q[0] ),
    .Y(_1624_));
 sky130_fd_sc_hd__a2111oi_1 _3649_ (.A1(_1619_),
    .A2(_1620_),
    .B1(_1622_),
    .C1(_1623_),
    .D1(_1624_),
    .Y(_1625_));
 sky130_fd_sc_hd__a32o_1 _3650_ (.A1(_1614_),
    .A2(_1617_),
    .A3(_1625_),
    .B1(_1624_),
    .B2(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_full_o ),
    .X(_0295_));
 sky130_fd_sc_hd__inv_2 _3651_ (.A(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_req_q ),
    .Y(_1626_));
 sky130_fd_sc_hd__or2_1 _3652_ (.A(_1626_),
    .B(_1235_),
    .X(_1627_));
 sky130_fd_sc_hd__a2bb2o_1 _3653_ (.A1_N(_1267_),
    .A2_N(_1627_),
    .B1(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_first_q[0] ),
    .B2(_1626_),
    .X(_1628_));
 sky130_fd_sc_hd__a21o_1 _3654_ (.A1(_2049_),
    .A2(_2078_),
    .B1(_1587_),
    .X(_1629_));
 sky130_fd_sc_hd__o21a_1 _3655_ (.A1(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_req_q ),
    .A2(\usb2uart.u_usb_cdc.bulk_in_req ),
    .B1(_1629_),
    .X(_1630_));
 sky130_fd_sc_hd__mux2_1 _3656_ (.A0(_1267_),
    .A1(_1628_),
    .S(_1630_),
    .X(_1631_));
 sky130_fd_sc_hd__clkbuf_1 _3657_ (.A(_1631_),
    .X(_0296_));
 sky130_fd_sc_hd__and2_1 _3658_ (.A(_1267_),
    .B(_1221_),
    .X(_1632_));
 sky130_fd_sc_hd__nor2_1 _3659_ (.A(_1234_),
    .B(_1632_),
    .Y(_1633_));
 sky130_fd_sc_hd__mux2_1 _3660_ (.A0(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_first_q[1] ),
    .A1(_1633_),
    .S(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_req_q ),
    .X(_1634_));
 sky130_fd_sc_hd__mux2_1 _3661_ (.A0(_1260_),
    .A1(_1634_),
    .S(_1630_),
    .X(_1635_));
 sky130_fd_sc_hd__clkbuf_1 _3662_ (.A(_1635_),
    .X(_0297_));
 sky130_fd_sc_hd__and3_1 _3663_ (.A(_1267_),
    .B(_1269_),
    .C(_1227_),
    .X(_1636_));
 sky130_fd_sc_hd__nor2_1 _3664_ (.A(_1265_),
    .B(_1632_),
    .Y(_1637_));
 sky130_fd_sc_hd__nor2_1 _3665_ (.A(_1636_),
    .B(_1637_),
    .Y(_1638_));
 sky130_fd_sc_hd__mux2_1 _3666_ (.A0(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_first_q[2] ),
    .A1(_1638_),
    .S(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_req_q ),
    .X(_1639_));
 sky130_fd_sc_hd__mux2_1 _3667_ (.A0(_1265_),
    .A1(_1639_),
    .S(_1630_),
    .X(_1640_));
 sky130_fd_sc_hd__clkbuf_1 _3668_ (.A(_1640_),
    .X(_0298_));
 sky130_fd_sc_hd__o21ai_1 _3669_ (.A1(_1627_),
    .A2(_1636_),
    .B1(_1630_),
    .Y(_1641_));
 sky130_fd_sc_hd__nor2_1 _3670_ (.A(_1626_),
    .B(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_first_qq[3] ),
    .Y(_1642_));
 sky130_fd_sc_hd__a22o_1 _3671_ (.A1(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_first_q[3] ),
    .A2(_1626_),
    .B1(_1636_),
    .B2(_1642_),
    .X(_1643_));
 sky130_fd_sc_hd__a22o_1 _3672_ (.A1(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_first_qq[3] ),
    .A2(_1641_),
    .B1(_1643_),
    .B2(_1630_),
    .X(_0299_));
 sky130_fd_sc_hd__and3_1 _3673_ (.A(_1626_),
    .B(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_state_q ),
    .C(_0779_),
    .X(_1644_));
 sky130_fd_sc_hd__and3_1 _3674_ (.A(\usb2uart.u_usb_cdc.in_data_ack ),
    .B(_1629_),
    .C(_1644_),
    .X(_1645_));
 sky130_fd_sc_hd__mux2_1 _3675_ (.A0(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_first_q[0] ),
    .A1(_1267_),
    .S(_1645_),
    .X(_1646_));
 sky130_fd_sc_hd__clkbuf_1 _3676_ (.A(_1646_),
    .X(_0300_));
 sky130_fd_sc_hd__mux2_1 _3677_ (.A0(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_first_q[1] ),
    .A1(_1260_),
    .S(_1645_),
    .X(_1647_));
 sky130_fd_sc_hd__clkbuf_1 _3678_ (.A(_1647_),
    .X(_0301_));
 sky130_fd_sc_hd__mux2_1 _3679_ (.A0(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_first_q[2] ),
    .A1(_1265_),
    .S(_1645_),
    .X(_1648_));
 sky130_fd_sc_hd__clkbuf_1 _3680_ (.A(_1648_),
    .X(_0302_));
 sky130_fd_sc_hd__mux2_1 _3681_ (.A0(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_first_q[3] ),
    .A1(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_first_qq[3] ),
    .S(_1645_),
    .X(_1649_));
 sky130_fd_sc_hd__clkbuf_1 _3682_ (.A(_1649_),
    .X(_0303_));
 sky130_fd_sc_hd__or3_1 _3683_ (.A(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_first_q[0] ),
    .B(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_first_q[1] ),
    .C(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_first_q[2] ),
    .X(_1650_));
 sky130_fd_sc_hd__nor2_1 _3684_ (.A(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_first_q[3] ),
    .B(_1650_),
    .Y(_1651_));
 sky130_fd_sc_hd__nor2_1 _3685_ (.A(_1591_),
    .B(_1651_),
    .Y(_1652_));
 sky130_fd_sc_hd__a21o_1 _3686_ (.A1(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_last_q[0] ),
    .A2(_1651_),
    .B1(_1652_),
    .X(_1653_));
 sky130_fd_sc_hd__nor2_1 _3687_ (.A(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_first_q[2] ),
    .B(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_first_q[3] ),
    .Y(_1654_));
 sky130_fd_sc_hd__or3_1 _3688_ (.A(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_first_q[0] ),
    .B(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_first_q[1] ),
    .C(_1654_),
    .X(_1655_));
 sky130_fd_sc_hd__xnor2_1 _3689_ (.A(_1592_),
    .B(_1655_),
    .Y(_1656_));
 sky130_fd_sc_hd__nand2_1 _3690_ (.A(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_first_q[0] ),
    .B(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_first_q[1] ),
    .Y(_1657_));
 sky130_fd_sc_hd__a21oi_1 _3691_ (.A1(_1655_),
    .A2(_1657_),
    .B1(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_last_q[1] ),
    .Y(_1658_));
 sky130_fd_sc_hd__xnor2_1 _3692_ (.A(_1588_),
    .B(_1650_),
    .Y(_1659_));
 sky130_fd_sc_hd__a31o_1 _3693_ (.A1(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_last_q[1] ),
    .A2(_1655_),
    .A3(_1657_),
    .B1(_1659_),
    .X(_1660_));
 sky130_fd_sc_hd__or4_2 _3694_ (.A(_1653_),
    .B(_1656_),
    .C(_1658_),
    .D(_1660_),
    .X(_1661_));
 sky130_fd_sc_hd__a21bo_1 _3695_ (.A1(\usb2uart.u_uart.uart_rx_inst.m_axis_tvalid_reg ),
    .A2(_1661_),
    .B1_N(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.delay_in_cnt_q[1] ),
    .X(_1662_));
 sky130_fd_sc_hd__nand2_1 _3696_ (.A(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.delay_in_cnt_q[0] ),
    .B(_1662_),
    .Y(_0304_));
 sky130_fd_sc_hd__and3_1 _3697_ (.A(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.delay_in_cnt_q[1] ),
    .B(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.delay_in_cnt_q[0] ),
    .C(_1661_),
    .X(_1663_));
 sky130_fd_sc_hd__and2_1 _3698_ (.A(\usb2uart.u_uart.uart_rx_inst.m_axis_tvalid_reg ),
    .B(_1663_),
    .X(_1664_));
 sky130_fd_sc_hd__buf_2 _3699_ (.A(_1664_),
    .X(_1665_));
 sky130_fd_sc_hd__clkbuf_4 _3700_ (.A(_1665_),
    .X(_1666_));
 sky130_fd_sc_hd__o21ba_1 _3701_ (.A1(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.delay_in_cnt_q[1] ),
    .A2(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.delay_in_cnt_q[0] ),
    .B1_N(_1666_),
    .X(_0305_));
 sky130_fd_sc_hd__or3_1 _3702_ (.A(\usb2uart.u_uart.uart_tx_inst.bit_cnt[3] ),
    .B(\usb2uart.u_uart.uart_tx_inst.bit_cnt[2] ),
    .C(\usb2uart.u_uart.uart_tx_inst.bit_cnt[1] ),
    .X(_1667_));
 sky130_fd_sc_hd__nor2_1 _3703_ (.A(\usb2uart.u_uart.uart_tx_inst.bit_cnt[0] ),
    .B(_1667_),
    .Y(_1668_));
 sky130_fd_sc_hd__buf_2 _3704_ (.A(_1668_),
    .X(_1669_));
 sky130_fd_sc_hd__buf_4 _3705_ (.A(_1594_),
    .X(_1670_));
 sky130_fd_sc_hd__mux2_1 _3706_ (.A0(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[16] ),
    .A1(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[24] ),
    .S(_1670_),
    .X(_1671_));
 sky130_fd_sc_hd__mux2_1 _3707_ (.A0(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[0] ),
    .A1(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[8] ),
    .S(_1594_),
    .X(_1672_));
 sky130_fd_sc_hd__and2b_1 _3708_ (.A_N(_1604_),
    .B(_1672_),
    .X(_1673_));
 sky130_fd_sc_hd__a211o_1 _3709_ (.A1(_1605_),
    .A2(_1671_),
    .B1(_1673_),
    .C1(_1609_),
    .X(_1674_));
 sky130_fd_sc_hd__buf_4 _3710_ (.A(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_first_q[0] ),
    .X(_1675_));
 sky130_fd_sc_hd__mux2_1 _3711_ (.A0(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[32] ),
    .A1(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[40] ),
    .S(_1675_),
    .X(_1676_));
 sky130_fd_sc_hd__and2b_1 _3712_ (.A_N(_1598_),
    .B(_1676_),
    .X(_1677_));
 sky130_fd_sc_hd__buf_2 _3713_ (.A(_1598_),
    .X(_1678_));
 sky130_fd_sc_hd__mux2_1 _3714_ (.A0(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[48] ),
    .A1(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[56] ),
    .S(_1675_),
    .X(_1679_));
 sky130_fd_sc_hd__and2_1 _3715_ (.A(_1678_),
    .B(_1679_),
    .X(_1680_));
 sky130_fd_sc_hd__o31a_1 _3716_ (.A1(_1610_),
    .A2(_1677_),
    .A3(_1680_),
    .B1(_1611_),
    .X(_1681_));
 sky130_fd_sc_hd__inv_2 _3717_ (.A(\usb2uart.u_uart.uart_tx_inst.bit_cnt[0] ),
    .Y(_1682_));
 sky130_fd_sc_hd__nor3_2 _3718_ (.A(\usb2uart.u_uart.uart_tx_inst.bit_cnt[3] ),
    .B(\usb2uart.u_uart.uart_tx_inst.bit_cnt[2] ),
    .C(\usb2uart.u_uart.uart_tx_inst.bit_cnt[1] ),
    .Y(_1683_));
 sky130_fd_sc_hd__nand2_4 _3719_ (.A(_1682_),
    .B(_1683_),
    .Y(_1684_));
 sky130_fd_sc_hd__a221o_1 _3720_ (.A1(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[64] ),
    .A2(_1602_),
    .B1(_1674_),
    .B2(_1681_),
    .C1(_1684_),
    .X(_1685_));
 sky130_fd_sc_hd__o21a_1 _3721_ (.A1(\usb2uart.u_uart.uart_tx_inst.data_reg[1] ),
    .A2(_1669_),
    .B1(_1685_),
    .X(_1686_));
 sky130_fd_sc_hd__or4_2 _3722_ (.A(\usb2uart.u_uart.uart_tx_inst.prescale_reg[3] ),
    .B(\usb2uart.u_uart.uart_tx_inst.prescale_reg[2] ),
    .C(\usb2uart.u_uart.uart_tx_inst.prescale_reg[1] ),
    .D(\usb2uart.u_uart.uart_tx_inst.prescale_reg[0] ),
    .X(_1687_));
 sky130_fd_sc_hd__or4_2 _3723_ (.A(\usb2uart.u_uart.uart_tx_inst.prescale_reg[6] ),
    .B(\usb2uart.u_uart.uart_tx_inst.prescale_reg[5] ),
    .C(\usb2uart.u_uart.uart_tx_inst.prescale_reg[4] ),
    .D(_1687_),
    .X(_1688_));
 sky130_fd_sc_hd__or2_1 _3724_ (.A(\usb2uart.u_uart.uart_tx_inst.prescale_reg[8] ),
    .B(\usb2uart.u_uart.uart_tx_inst.prescale_reg[7] ),
    .X(_1689_));
 sky130_fd_sc_hd__or4_2 _3725_ (.A(\usb2uart.u_uart.uart_tx_inst.prescale_reg[10] ),
    .B(\usb2uart.u_uart.uart_tx_inst.prescale_reg[9] ),
    .C(_1688_),
    .D(_1689_),
    .X(_1690_));
 sky130_fd_sc_hd__or4_2 _3726_ (.A(\usb2uart.u_uart.uart_tx_inst.prescale_reg[13] ),
    .B(\usb2uart.u_uart.uart_tx_inst.prescale_reg[12] ),
    .C(\usb2uart.u_uart.uart_tx_inst.prescale_reg[11] ),
    .D(_1690_),
    .X(_1691_));
 sky130_fd_sc_hd__or4_1 _3727_ (.A(\usb2uart.u_uart.uart_tx_inst.prescale_reg[16] ),
    .B(\usb2uart.u_uart.uart_tx_inst.prescale_reg[15] ),
    .C(\usb2uart.u_uart.uart_tx_inst.prescale_reg[14] ),
    .D(_1691_),
    .X(_1692_));
 sky130_fd_sc_hd__or2_1 _3728_ (.A(\usb2uart.u_uart.uart_tx_inst.prescale_reg[17] ),
    .B(_1692_),
    .X(_1693_));
 sky130_fd_sc_hd__nor2_2 _3729_ (.A(\usb2uart.u_uart.uart_tx_inst.prescale_reg[18] ),
    .B(_1693_),
    .Y(_1694_));
 sky130_fd_sc_hd__a31o_1 _3730_ (.A1(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.delay_out_cnt_q[1] ),
    .A2(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.delay_out_cnt_q[0] ),
    .A3(_1578_),
    .B1(_1684_),
    .X(_1695_));
 sky130_fd_sc_hd__nand2_1 _3731_ (.A(_1694_),
    .B(_1695_),
    .Y(_1696_));
 sky130_fd_sc_hd__or2_1 _3732_ (.A(\usb2uart.u_uart.uart_tx_inst.prescale_reg[18] ),
    .B(_1693_),
    .X(_1697_));
 sky130_fd_sc_hd__or2_2 _3733_ (.A(_1697_),
    .B(_1695_),
    .X(_1698_));
 sky130_fd_sc_hd__o21ai_1 _3734_ (.A1(_1682_),
    .A2(_1667_),
    .B1(_1694_),
    .Y(_1699_));
 sky130_fd_sc_hd__o21ai_1 _3735_ (.A1(\usb2uart.u_uart.uart_tx_inst.prescale_reg[0] ),
    .A2(_1694_),
    .B1(_1699_),
    .Y(_1700_));
 sky130_fd_sc_hd__nand2_1 _3736_ (.A(_1698_),
    .B(_1700_),
    .Y(_1701_));
 sky130_fd_sc_hd__or3_1 _3737_ (.A(net4),
    .B(_1696_),
    .C(_1701_),
    .X(_1702_));
 sky130_fd_sc_hd__clkbuf_4 _3738_ (.A(_1702_),
    .X(_1703_));
 sky130_fd_sc_hd__mux2_1 _3739_ (.A0(_1686_),
    .A1(\usb2uart.u_uart.uart_tx_inst.data_reg[0] ),
    .S(_1703_),
    .X(_1704_));
 sky130_fd_sc_hd__clkbuf_1 _3740_ (.A(_1704_),
    .X(_0306_));
 sky130_fd_sc_hd__mux2_1 _3741_ (.A0(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[17] ),
    .A1(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[25] ),
    .S(_1670_),
    .X(_1705_));
 sky130_fd_sc_hd__mux2_1 _3742_ (.A0(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[1] ),
    .A1(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[9] ),
    .S(_1594_),
    .X(_1706_));
 sky130_fd_sc_hd__and2b_1 _3743_ (.A_N(_1604_),
    .B(_1706_),
    .X(_1707_));
 sky130_fd_sc_hd__a211o_1 _3744_ (.A1(_1605_),
    .A2(_1705_),
    .B1(_1707_),
    .C1(_1609_),
    .X(_1708_));
 sky130_fd_sc_hd__or2b_1 _3745_ (.A(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[41] ),
    .B_N(_1595_),
    .X(_1709_));
 sky130_fd_sc_hd__o21ba_1 _3746_ (.A1(_1595_),
    .A2(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[33] ),
    .B1_N(_1678_),
    .X(_1710_));
 sky130_fd_sc_hd__mux2_1 _3747_ (.A0(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[49] ),
    .A1(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[57] ),
    .S(_1670_),
    .X(_1711_));
 sky130_fd_sc_hd__a221o_1 _3748_ (.A1(_1709_),
    .A2(_1710_),
    .B1(_1711_),
    .B2(_1604_),
    .C1(_1610_),
    .X(_1712_));
 sky130_fd_sc_hd__a21o_1 _3749_ (.A1(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[65] ),
    .A2(_1602_),
    .B1(_1684_),
    .X(_1713_));
 sky130_fd_sc_hd__a31o_1 _3750_ (.A1(_1611_),
    .A2(_1708_),
    .A3(_1712_),
    .B1(_1713_),
    .X(_1714_));
 sky130_fd_sc_hd__o21a_1 _3751_ (.A1(\usb2uart.u_uart.uart_tx_inst.data_reg[2] ),
    .A2(_1669_),
    .B1(_1714_),
    .X(_1715_));
 sky130_fd_sc_hd__mux2_1 _3752_ (.A0(_1715_),
    .A1(\usb2uart.u_uart.uart_tx_inst.data_reg[1] ),
    .S(_1703_),
    .X(_1716_));
 sky130_fd_sc_hd__clkbuf_1 _3753_ (.A(_1716_),
    .X(_0307_));
 sky130_fd_sc_hd__mux2_1 _3754_ (.A0(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[18] ),
    .A1(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[26] ),
    .S(_1670_),
    .X(_1717_));
 sky130_fd_sc_hd__mux2_1 _3755_ (.A0(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[2] ),
    .A1(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[10] ),
    .S(_1594_),
    .X(_1718_));
 sky130_fd_sc_hd__and2b_1 _3756_ (.A_N(_1678_),
    .B(_1718_),
    .X(_1719_));
 sky130_fd_sc_hd__a211o_1 _3757_ (.A1(_1605_),
    .A2(_1717_),
    .B1(_1719_),
    .C1(_1609_),
    .X(_1720_));
 sky130_fd_sc_hd__mux2_1 _3758_ (.A0(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[34] ),
    .A1(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[42] ),
    .S(_1675_),
    .X(_1721_));
 sky130_fd_sc_hd__and2b_1 _3759_ (.A_N(_1598_),
    .B(_1721_),
    .X(_1722_));
 sky130_fd_sc_hd__mux2_1 _3760_ (.A0(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[50] ),
    .A1(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[58] ),
    .S(_1675_),
    .X(_1723_));
 sky130_fd_sc_hd__and2_1 _3761_ (.A(_1678_),
    .B(_1723_),
    .X(_1724_));
 sky130_fd_sc_hd__o31a_1 _3762_ (.A1(_1610_),
    .A2(_1722_),
    .A3(_1724_),
    .B1(_1611_),
    .X(_1725_));
 sky130_fd_sc_hd__a221o_1 _3763_ (.A1(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[66] ),
    .A2(_1602_),
    .B1(_1720_),
    .B2(_1725_),
    .C1(_1684_),
    .X(_1726_));
 sky130_fd_sc_hd__o21a_1 _3764_ (.A1(\usb2uart.u_uart.uart_tx_inst.data_reg[3] ),
    .A2(_1669_),
    .B1(_1726_),
    .X(_1727_));
 sky130_fd_sc_hd__mux2_1 _3765_ (.A0(_1727_),
    .A1(\usb2uart.u_uart.uart_tx_inst.data_reg[2] ),
    .S(_1703_),
    .X(_1728_));
 sky130_fd_sc_hd__clkbuf_1 _3766_ (.A(_1728_),
    .X(_0308_));
 sky130_fd_sc_hd__mux2_1 _3767_ (.A0(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[19] ),
    .A1(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[27] ),
    .S(_1670_),
    .X(_1729_));
 sky130_fd_sc_hd__mux2_1 _3768_ (.A0(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[3] ),
    .A1(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[11] ),
    .S(_1594_),
    .X(_1730_));
 sky130_fd_sc_hd__and2b_1 _3769_ (.A_N(_1678_),
    .B(_1730_),
    .X(_1731_));
 sky130_fd_sc_hd__a211o_1 _3770_ (.A1(_1605_),
    .A2(_1729_),
    .B1(_1731_),
    .C1(_1609_),
    .X(_1732_));
 sky130_fd_sc_hd__mux2_1 _3771_ (.A0(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[35] ),
    .A1(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[43] ),
    .S(_1675_),
    .X(_1733_));
 sky130_fd_sc_hd__and2b_1 _3772_ (.A_N(_1598_),
    .B(_1733_),
    .X(_1734_));
 sky130_fd_sc_hd__mux2_1 _3773_ (.A0(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[51] ),
    .A1(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[59] ),
    .S(_1675_),
    .X(_1735_));
 sky130_fd_sc_hd__and2_1 _3774_ (.A(_1678_),
    .B(_1735_),
    .X(_1736_));
 sky130_fd_sc_hd__o31a_1 _3775_ (.A1(_1610_),
    .A2(_1734_),
    .A3(_1736_),
    .B1(_1611_),
    .X(_1737_));
 sky130_fd_sc_hd__a221o_1 _3776_ (.A1(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[67] ),
    .A2(_1602_),
    .B1(_1732_),
    .B2(_1737_),
    .C1(_1684_),
    .X(_1738_));
 sky130_fd_sc_hd__o21a_1 _3777_ (.A1(\usb2uart.u_uart.uart_tx_inst.data_reg[4] ),
    .A2(_1669_),
    .B1(_1738_),
    .X(_1739_));
 sky130_fd_sc_hd__mux2_1 _3778_ (.A0(_1739_),
    .A1(\usb2uart.u_uart.uart_tx_inst.data_reg[3] ),
    .S(_1703_),
    .X(_1740_));
 sky130_fd_sc_hd__clkbuf_1 _3779_ (.A(_1740_),
    .X(_0309_));
 sky130_fd_sc_hd__mux2_1 _3780_ (.A0(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[20] ),
    .A1(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[28] ),
    .S(_1670_),
    .X(_1741_));
 sky130_fd_sc_hd__mux2_1 _3781_ (.A0(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[4] ),
    .A1(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[12] ),
    .S(_1594_),
    .X(_1742_));
 sky130_fd_sc_hd__and2b_1 _3782_ (.A_N(_1604_),
    .B(_1742_),
    .X(_1743_));
 sky130_fd_sc_hd__a211o_1 _3783_ (.A1(_1605_),
    .A2(_1741_),
    .B1(_1743_),
    .C1(_1609_),
    .X(_1744_));
 sky130_fd_sc_hd__or2b_1 _3784_ (.A(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[44] ),
    .B_N(_1595_),
    .X(_1745_));
 sky130_fd_sc_hd__o21ba_1 _3785_ (.A1(_1595_),
    .A2(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[36] ),
    .B1_N(_1598_),
    .X(_1746_));
 sky130_fd_sc_hd__mux2_1 _3786_ (.A0(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[52] ),
    .A1(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[60] ),
    .S(_1670_),
    .X(_1747_));
 sky130_fd_sc_hd__a221o_1 _3787_ (.A1(_1745_),
    .A2(_1746_),
    .B1(_1747_),
    .B2(_1604_),
    .C1(_1610_),
    .X(_1748_));
 sky130_fd_sc_hd__a21o_1 _3788_ (.A1(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[68] ),
    .A2(_1602_),
    .B1(_1684_),
    .X(_1749_));
 sky130_fd_sc_hd__a31o_1 _3789_ (.A1(_1611_),
    .A2(_1744_),
    .A3(_1748_),
    .B1(_1749_),
    .X(_1750_));
 sky130_fd_sc_hd__o21a_1 _3790_ (.A1(\usb2uart.u_uart.uart_tx_inst.data_reg[5] ),
    .A2(_1669_),
    .B1(_1750_),
    .X(_1751_));
 sky130_fd_sc_hd__mux2_1 _3791_ (.A0(_1751_),
    .A1(\usb2uart.u_uart.uart_tx_inst.data_reg[4] ),
    .S(_1703_),
    .X(_1752_));
 sky130_fd_sc_hd__clkbuf_1 _3792_ (.A(_1752_),
    .X(_0310_));
 sky130_fd_sc_hd__mux2_1 _3793_ (.A0(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[21] ),
    .A1(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[29] ),
    .S(_1594_),
    .X(_1753_));
 sky130_fd_sc_hd__mux2_1 _3794_ (.A0(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[5] ),
    .A1(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[13] ),
    .S(_1675_),
    .X(_1754_));
 sky130_fd_sc_hd__and2b_1 _3795_ (.A_N(_1678_),
    .B(_1754_),
    .X(_1755_));
 sky130_fd_sc_hd__a211o_1 _3796_ (.A1(_1604_),
    .A2(_1753_),
    .B1(_1755_),
    .C1(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_first_q[2] ),
    .X(_1756_));
 sky130_fd_sc_hd__mux2_1 _3797_ (.A0(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[37] ),
    .A1(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[45] ),
    .S(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_first_q[0] ),
    .X(_1757_));
 sky130_fd_sc_hd__and2b_1 _3798_ (.A_N(_1598_),
    .B(_1757_),
    .X(_1758_));
 sky130_fd_sc_hd__mux2_1 _3799_ (.A0(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[53] ),
    .A1(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[61] ),
    .S(_1675_),
    .X(_1759_));
 sky130_fd_sc_hd__and2_1 _3800_ (.A(_1678_),
    .B(_1759_),
    .X(_1760_));
 sky130_fd_sc_hd__o31a_1 _3801_ (.A1(_1610_),
    .A2(_1758_),
    .A3(_1760_),
    .B1(_1611_),
    .X(_1761_));
 sky130_fd_sc_hd__a221o_1 _3802_ (.A1(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[69] ),
    .A2(_1602_),
    .B1(_1756_),
    .B2(_1761_),
    .C1(_1684_),
    .X(_1762_));
 sky130_fd_sc_hd__o21a_1 _3803_ (.A1(\usb2uart.u_uart.uart_tx_inst.data_reg[6] ),
    .A2(_1669_),
    .B1(_1762_),
    .X(_1763_));
 sky130_fd_sc_hd__mux2_1 _3804_ (.A0(_1763_),
    .A1(\usb2uart.u_uart.uart_tx_inst.data_reg[5] ),
    .S(_1703_),
    .X(_1764_));
 sky130_fd_sc_hd__clkbuf_1 _3805_ (.A(_1764_),
    .X(_0311_));
 sky130_fd_sc_hd__mux2_1 _3806_ (.A0(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[22] ),
    .A1(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[30] ),
    .S(_1594_),
    .X(_1765_));
 sky130_fd_sc_hd__mux2_1 _3807_ (.A0(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[6] ),
    .A1(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[14] ),
    .S(_1675_),
    .X(_1766_));
 sky130_fd_sc_hd__and2b_1 _3808_ (.A_N(_1678_),
    .B(_1766_),
    .X(_1767_));
 sky130_fd_sc_hd__a211o_1 _3809_ (.A1(_1604_),
    .A2(_1765_),
    .B1(_1767_),
    .C1(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_first_q[2] ),
    .X(_1768_));
 sky130_fd_sc_hd__mux2_1 _3810_ (.A0(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[38] ),
    .A1(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[46] ),
    .S(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_first_q[0] ),
    .X(_1769_));
 sky130_fd_sc_hd__and2b_1 _3811_ (.A_N(_1598_),
    .B(_1769_),
    .X(_1770_));
 sky130_fd_sc_hd__mux2_1 _3812_ (.A0(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[54] ),
    .A1(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[62] ),
    .S(_1675_),
    .X(_1771_));
 sky130_fd_sc_hd__and2_1 _3813_ (.A(_1678_),
    .B(_1771_),
    .X(_1772_));
 sky130_fd_sc_hd__o31a_1 _3814_ (.A1(_1610_),
    .A2(_1770_),
    .A3(_1772_),
    .B1(_1611_),
    .X(_1773_));
 sky130_fd_sc_hd__a221o_1 _3815_ (.A1(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[70] ),
    .A2(_1602_),
    .B1(_1768_),
    .B2(_1773_),
    .C1(_1684_),
    .X(_1774_));
 sky130_fd_sc_hd__o21a_1 _3816_ (.A1(\usb2uart.u_uart.uart_tx_inst.data_reg[7] ),
    .A2(_1669_),
    .B1(_1774_),
    .X(_1775_));
 sky130_fd_sc_hd__mux2_1 _3817_ (.A0(_1775_),
    .A1(\usb2uart.u_uart.uart_tx_inst.data_reg[6] ),
    .S(_1703_),
    .X(_1776_));
 sky130_fd_sc_hd__clkbuf_1 _3818_ (.A(_1776_),
    .X(_0312_));
 sky130_fd_sc_hd__mux2_1 _3819_ (.A0(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[23] ),
    .A1(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[31] ),
    .S(_1670_),
    .X(_1777_));
 sky130_fd_sc_hd__mux2_1 _3820_ (.A0(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[7] ),
    .A1(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[15] ),
    .S(_1594_),
    .X(_1778_));
 sky130_fd_sc_hd__and2b_1 _3821_ (.A_N(_1604_),
    .B(_1778_),
    .X(_1779_));
 sky130_fd_sc_hd__a211o_1 _3822_ (.A1(_1605_),
    .A2(_1777_),
    .B1(_1779_),
    .C1(_1609_),
    .X(_1780_));
 sky130_fd_sc_hd__or2b_1 _3823_ (.A(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[47] ),
    .B_N(_1595_),
    .X(_1781_));
 sky130_fd_sc_hd__o21ba_1 _3824_ (.A1(_1670_),
    .A2(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[39] ),
    .B1_N(_1598_),
    .X(_1782_));
 sky130_fd_sc_hd__mux2_1 _3825_ (.A0(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[55] ),
    .A1(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[63] ),
    .S(_1670_),
    .X(_1783_));
 sky130_fd_sc_hd__a221o_1 _3826_ (.A1(_1781_),
    .A2(_1782_),
    .B1(_1783_),
    .B2(_1604_),
    .C1(_1610_),
    .X(_1784_));
 sky130_fd_sc_hd__a21o_1 _3827_ (.A1(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[71] ),
    .A2(_1602_),
    .B1(_1684_),
    .X(_1785_));
 sky130_fd_sc_hd__a31o_1 _3828_ (.A1(_1611_),
    .A2(_1780_),
    .A3(_1784_),
    .B1(_1785_),
    .X(_1786_));
 sky130_fd_sc_hd__o21a_1 _3829_ (.A1(\usb2uart.u_uart.uart_tx_inst.data_reg[8] ),
    .A2(_1668_),
    .B1(_1786_),
    .X(_1787_));
 sky130_fd_sc_hd__mux2_1 _3830_ (.A0(_1787_),
    .A1(\usb2uart.u_uart.uart_tx_inst.data_reg[7] ),
    .S(_1703_),
    .X(_1788_));
 sky130_fd_sc_hd__clkbuf_1 _3831_ (.A(_1788_),
    .X(_0313_));
 sky130_fd_sc_hd__mux2_1 _3832_ (.A0(_1669_),
    .A1(\usb2uart.u_uart.uart_tx_inst.data_reg[8] ),
    .S(_1703_),
    .X(_1789_));
 sky130_fd_sc_hd__clkbuf_1 _3833_ (.A(_1789_),
    .X(_0314_));
 sky130_fd_sc_hd__or3_4 _3834_ (.A(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_last_q[1] ),
    .B(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_last_q[2] ),
    .C(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_last_q[3] ),
    .X(_1790_));
 sky130_fd_sc_hd__or3b_1 _3835_ (.A(_1790_),
    .B(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_last_q[0] ),
    .C_N(_1665_),
    .X(_1791_));
 sky130_fd_sc_hd__clkbuf_4 _3836_ (.A(_1791_),
    .X(_1792_));
 sky130_fd_sc_hd__mux2_1 _3837_ (.A0(\usb2uart.u_uart.uart_rx_inst.m_axis_tdata_reg[0] ),
    .A1(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[0] ),
    .S(_1792_),
    .X(_1793_));
 sky130_fd_sc_hd__clkbuf_1 _3838_ (.A(_1793_),
    .X(_0315_));
 sky130_fd_sc_hd__mux2_1 _3839_ (.A0(\usb2uart.u_uart.uart_rx_inst.m_axis_tdata_reg[1] ),
    .A1(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[1] ),
    .S(_1792_),
    .X(_1794_));
 sky130_fd_sc_hd__clkbuf_1 _3840_ (.A(_1794_),
    .X(_0316_));
 sky130_fd_sc_hd__mux2_1 _3841_ (.A0(\usb2uart.u_uart.uart_rx_inst.m_axis_tdata_reg[2] ),
    .A1(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[2] ),
    .S(_1792_),
    .X(_1795_));
 sky130_fd_sc_hd__clkbuf_1 _3842_ (.A(_1795_),
    .X(_0317_));
 sky130_fd_sc_hd__mux2_1 _3843_ (.A0(\usb2uart.u_uart.uart_rx_inst.m_axis_tdata_reg[3] ),
    .A1(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[3] ),
    .S(_1792_),
    .X(_1796_));
 sky130_fd_sc_hd__clkbuf_1 _3844_ (.A(_1796_),
    .X(_0318_));
 sky130_fd_sc_hd__mux2_1 _3845_ (.A0(\usb2uart.u_uart.uart_rx_inst.m_axis_tdata_reg[4] ),
    .A1(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[4] ),
    .S(_1792_),
    .X(_1797_));
 sky130_fd_sc_hd__clkbuf_1 _3846_ (.A(_1797_),
    .X(_0319_));
 sky130_fd_sc_hd__mux2_1 _3847_ (.A0(\usb2uart.u_uart.uart_rx_inst.m_axis_tdata_reg[5] ),
    .A1(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[5] ),
    .S(_1792_),
    .X(_1798_));
 sky130_fd_sc_hd__clkbuf_1 _3848_ (.A(_1798_),
    .X(_0320_));
 sky130_fd_sc_hd__mux2_1 _3849_ (.A0(\usb2uart.u_uart.uart_rx_inst.m_axis_tdata_reg[6] ),
    .A1(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[6] ),
    .S(_1792_),
    .X(_1799_));
 sky130_fd_sc_hd__clkbuf_1 _3850_ (.A(_1799_),
    .X(_0321_));
 sky130_fd_sc_hd__mux2_1 _3851_ (.A0(\usb2uart.u_uart.uart_rx_inst.m_axis_tdata_reg[7] ),
    .A1(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[7] ),
    .S(_1792_),
    .X(_1800_));
 sky130_fd_sc_hd__clkbuf_1 _3852_ (.A(_1800_),
    .X(_0322_));
 sky130_fd_sc_hd__nand2_1 _3853_ (.A(_1582_),
    .B(_1665_),
    .Y(_1801_));
 sky130_fd_sc_hd__or2_1 _3854_ (.A(_1790_),
    .B(_1801_),
    .X(_1802_));
 sky130_fd_sc_hd__buf_2 _3855_ (.A(_1802_),
    .X(_1803_));
 sky130_fd_sc_hd__or2_2 _3856_ (.A(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_last_q[0] ),
    .B(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_last_q[1] ),
    .X(_1804_));
 sky130_fd_sc_hd__nor2_1 _3857_ (.A(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_last_q[2] ),
    .B(_1804_),
    .Y(_1805_));
 sky130_fd_sc_hd__clkbuf_4 _3858_ (.A(_1805_),
    .X(_1806_));
 sky130_fd_sc_hd__nand2_1 _3859_ (.A(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_last_q[2] ),
    .B(_1804_),
    .Y(_1807_));
 sky130_fd_sc_hd__nand3b_2 _3860_ (.A_N(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_last_q[3] ),
    .B(_1665_),
    .C(_1807_),
    .Y(_1808_));
 sky130_fd_sc_hd__nor2_4 _3861_ (.A(_1806_),
    .B(_1808_),
    .Y(_1809_));
 sky130_fd_sc_hd__buf_2 _3862_ (.A(_1582_),
    .X(_1810_));
 sky130_fd_sc_hd__and3b_1 _3863_ (.A_N(_1589_),
    .B(_1810_),
    .C(\usb2uart.u_uart.uart_rx_inst.m_axis_tdata_reg[0] ),
    .X(_1811_));
 sky130_fd_sc_hd__a22o_1 _3864_ (.A1(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[8] ),
    .A2(_1803_),
    .B1(_1809_),
    .B2(_1811_),
    .X(_0323_));
 sky130_fd_sc_hd__and3b_1 _3865_ (.A_N(_1589_),
    .B(_1582_),
    .C(\usb2uart.u_uart.uart_rx_inst.m_axis_tdata_reg[1] ),
    .X(_1812_));
 sky130_fd_sc_hd__a22o_1 _3866_ (.A1(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[9] ),
    .A2(_1803_),
    .B1(_1809_),
    .B2(_1812_),
    .X(_0324_));
 sky130_fd_sc_hd__and3b_1 _3867_ (.A_N(_1589_),
    .B(_1582_),
    .C(\usb2uart.u_uart.uart_rx_inst.m_axis_tdata_reg[2] ),
    .X(_1813_));
 sky130_fd_sc_hd__a22o_1 _3868_ (.A1(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[10] ),
    .A2(_1803_),
    .B1(_1809_),
    .B2(_1813_),
    .X(_0325_));
 sky130_fd_sc_hd__and3b_1 _3869_ (.A_N(_1589_),
    .B(_1582_),
    .C(\usb2uart.u_uart.uart_rx_inst.m_axis_tdata_reg[3] ),
    .X(_1814_));
 sky130_fd_sc_hd__a22o_1 _3870_ (.A1(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[11] ),
    .A2(_1803_),
    .B1(_1809_),
    .B2(_1814_),
    .X(_0326_));
 sky130_fd_sc_hd__and3b_1 _3871_ (.A_N(_1589_),
    .B(_1582_),
    .C(\usb2uart.u_uart.uart_rx_inst.m_axis_tdata_reg[4] ),
    .X(_1815_));
 sky130_fd_sc_hd__a22o_1 _3872_ (.A1(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[12] ),
    .A2(_1803_),
    .B1(_1809_),
    .B2(_1815_),
    .X(_0327_));
 sky130_fd_sc_hd__and3b_1 _3873_ (.A_N(_1589_),
    .B(_1582_),
    .C(\usb2uart.u_uart.uart_rx_inst.m_axis_tdata_reg[5] ),
    .X(_1816_));
 sky130_fd_sc_hd__a22o_1 _3874_ (.A1(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[13] ),
    .A2(_1803_),
    .B1(_1809_),
    .B2(_1816_),
    .X(_0328_));
 sky130_fd_sc_hd__and3b_1 _3875_ (.A_N(_1589_),
    .B(_1582_),
    .C(\usb2uart.u_uart.uart_rx_inst.m_axis_tdata_reg[6] ),
    .X(_1817_));
 sky130_fd_sc_hd__a22o_1 _3876_ (.A1(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[14] ),
    .A2(_1803_),
    .B1(_1809_),
    .B2(_1817_),
    .X(_0329_));
 sky130_fd_sc_hd__and2b_1 _3877_ (.A_N(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_last_q[1] ),
    .B(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_last_q[0] ),
    .X(_1818_));
 sky130_fd_sc_hd__a32o_1 _3878_ (.A1(\usb2uart.u_uart.uart_rx_inst.m_axis_tdata_reg[7] ),
    .A2(_1809_),
    .A3(_1818_),
    .B1(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[15] ),
    .B2(_1803_),
    .X(_0330_));
 sky130_fd_sc_hd__and2_1 _3879_ (.A(\usb2uart.u_uart.uart_rx_inst.m_axis_tdata_reg[0] ),
    .B(_1790_),
    .X(_1819_));
 sky130_fd_sc_hd__or3b_1 _3880_ (.A(_1808_),
    .B(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_last_q[0] ),
    .C_N(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_last_q[1] ),
    .X(_1820_));
 sky130_fd_sc_hd__clkbuf_4 _3881_ (.A(_1820_),
    .X(_1821_));
 sky130_fd_sc_hd__mux2_1 _3882_ (.A0(_1819_),
    .A1(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[16] ),
    .S(_1821_),
    .X(_1822_));
 sky130_fd_sc_hd__clkbuf_1 _3883_ (.A(_1822_),
    .X(_0331_));
 sky130_fd_sc_hd__and2_1 _3884_ (.A(\usb2uart.u_uart.uart_rx_inst.m_axis_tdata_reg[1] ),
    .B(_1790_),
    .X(_1823_));
 sky130_fd_sc_hd__mux2_1 _3885_ (.A0(_1823_),
    .A1(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[17] ),
    .S(_1821_),
    .X(_1824_));
 sky130_fd_sc_hd__clkbuf_1 _3886_ (.A(_1824_),
    .X(_0332_));
 sky130_fd_sc_hd__and2_1 _3887_ (.A(\usb2uart.u_uart.uart_rx_inst.m_axis_tdata_reg[2] ),
    .B(_1790_),
    .X(_1825_));
 sky130_fd_sc_hd__mux2_1 _3888_ (.A0(_1825_),
    .A1(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[18] ),
    .S(_1821_),
    .X(_1826_));
 sky130_fd_sc_hd__clkbuf_1 _3889_ (.A(_1826_),
    .X(_0333_));
 sky130_fd_sc_hd__and2_1 _3890_ (.A(\usb2uart.u_uart.uart_rx_inst.m_axis_tdata_reg[3] ),
    .B(_1790_),
    .X(_1827_));
 sky130_fd_sc_hd__mux2_1 _3891_ (.A0(_1827_),
    .A1(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[19] ),
    .S(_1821_),
    .X(_1828_));
 sky130_fd_sc_hd__clkbuf_1 _3892_ (.A(_1828_),
    .X(_0334_));
 sky130_fd_sc_hd__and2_1 _3893_ (.A(\usb2uart.u_uart.uart_rx_inst.m_axis_tdata_reg[4] ),
    .B(_1790_),
    .X(_1829_));
 sky130_fd_sc_hd__mux2_1 _3894_ (.A0(_1829_),
    .A1(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[20] ),
    .S(_1821_),
    .X(_1830_));
 sky130_fd_sc_hd__clkbuf_1 _3895_ (.A(_1830_),
    .X(_0335_));
 sky130_fd_sc_hd__and2_1 _3896_ (.A(\usb2uart.u_uart.uart_rx_inst.m_axis_tdata_reg[5] ),
    .B(_1790_),
    .X(_1831_));
 sky130_fd_sc_hd__mux2_1 _3897_ (.A0(_1831_),
    .A1(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[21] ),
    .S(_1821_),
    .X(_1832_));
 sky130_fd_sc_hd__clkbuf_1 _3898_ (.A(_1832_),
    .X(_0336_));
 sky130_fd_sc_hd__and2_1 _3899_ (.A(\usb2uart.u_uart.uart_rx_inst.m_axis_tdata_reg[6] ),
    .B(_1790_),
    .X(_1833_));
 sky130_fd_sc_hd__mux2_1 _3900_ (.A0(_1833_),
    .A1(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[22] ),
    .S(_1821_),
    .X(_1834_));
 sky130_fd_sc_hd__clkbuf_1 _3901_ (.A(_1834_),
    .X(_0337_));
 sky130_fd_sc_hd__and2_1 _3902_ (.A(\usb2uart.u_uart.uart_rx_inst.m_axis_tdata_reg[7] ),
    .B(_1790_),
    .X(_1835_));
 sky130_fd_sc_hd__mux2_1 _3903_ (.A0(_1835_),
    .A1(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[23] ),
    .S(_1821_),
    .X(_1836_));
 sky130_fd_sc_hd__clkbuf_1 _3904_ (.A(_1836_),
    .X(_0338_));
 sky130_fd_sc_hd__nand2_1 _3905_ (.A(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_last_q[0] ),
    .B(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_last_q[1] ),
    .Y(_1837_));
 sky130_fd_sc_hd__or2_1 _3906_ (.A(_1808_),
    .B(_1837_),
    .X(_1838_));
 sky130_fd_sc_hd__buf_4 _3907_ (.A(_1838_),
    .X(_1839_));
 sky130_fd_sc_hd__mux2_1 _3908_ (.A0(\usb2uart.u_uart.uart_rx_inst.m_axis_tdata_reg[0] ),
    .A1(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[24] ),
    .S(_1839_),
    .X(_1840_));
 sky130_fd_sc_hd__clkbuf_1 _3909_ (.A(_1840_),
    .X(_0339_));
 sky130_fd_sc_hd__mux2_1 _3910_ (.A0(\usb2uart.u_uart.uart_rx_inst.m_axis_tdata_reg[1] ),
    .A1(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[25] ),
    .S(_1839_),
    .X(_1841_));
 sky130_fd_sc_hd__clkbuf_1 _3911_ (.A(_1841_),
    .X(_0340_));
 sky130_fd_sc_hd__mux2_1 _3912_ (.A0(\usb2uart.u_uart.uart_rx_inst.m_axis_tdata_reg[2] ),
    .A1(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[26] ),
    .S(_1839_),
    .X(_1842_));
 sky130_fd_sc_hd__clkbuf_1 _3913_ (.A(_1842_),
    .X(_0341_));
 sky130_fd_sc_hd__mux2_1 _3914_ (.A0(\usb2uart.u_uart.uart_rx_inst.m_axis_tdata_reg[3] ),
    .A1(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[27] ),
    .S(_1839_),
    .X(_1843_));
 sky130_fd_sc_hd__clkbuf_1 _3915_ (.A(_1843_),
    .X(_0342_));
 sky130_fd_sc_hd__mux2_1 _3916_ (.A0(\usb2uart.u_uart.uart_rx_inst.m_axis_tdata_reg[4] ),
    .A1(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[28] ),
    .S(_1839_),
    .X(_1844_));
 sky130_fd_sc_hd__clkbuf_1 _3917_ (.A(_1844_),
    .X(_0343_));
 sky130_fd_sc_hd__mux2_1 _3918_ (.A0(\usb2uart.u_uart.uart_rx_inst.m_axis_tdata_reg[5] ),
    .A1(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[29] ),
    .S(_1839_),
    .X(_1845_));
 sky130_fd_sc_hd__clkbuf_1 _3919_ (.A(_1845_),
    .X(_0344_));
 sky130_fd_sc_hd__mux2_1 _3920_ (.A0(\usb2uart.u_uart.uart_rx_inst.m_axis_tdata_reg[6] ),
    .A1(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[30] ),
    .S(_1839_),
    .X(_1846_));
 sky130_fd_sc_hd__clkbuf_1 _3921_ (.A(_1846_),
    .X(_0345_));
 sky130_fd_sc_hd__mux2_1 _3922_ (.A0(\usb2uart.u_uart.uart_rx_inst.m_axis_tdata_reg[7] ),
    .A1(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[31] ),
    .S(_1839_),
    .X(_1847_));
 sky130_fd_sc_hd__clkbuf_1 _3923_ (.A(_1847_),
    .X(_0346_));
 sky130_fd_sc_hd__or3_1 _3924_ (.A(_1804_),
    .B(_1806_),
    .C(_1808_),
    .X(_1848_));
 sky130_fd_sc_hd__clkbuf_4 _3925_ (.A(_1848_),
    .X(_1849_));
 sky130_fd_sc_hd__mux2_1 _3926_ (.A0(_1819_),
    .A1(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[32] ),
    .S(_1849_),
    .X(_1850_));
 sky130_fd_sc_hd__clkbuf_1 _3927_ (.A(_1850_),
    .X(_0347_));
 sky130_fd_sc_hd__mux2_1 _3928_ (.A0(_1823_),
    .A1(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[33] ),
    .S(_1849_),
    .X(_1851_));
 sky130_fd_sc_hd__clkbuf_1 _3929_ (.A(_1851_),
    .X(_0348_));
 sky130_fd_sc_hd__mux2_1 _3930_ (.A0(_1825_),
    .A1(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[34] ),
    .S(_1849_),
    .X(_1852_));
 sky130_fd_sc_hd__clkbuf_1 _3931_ (.A(_1852_),
    .X(_0349_));
 sky130_fd_sc_hd__mux2_1 _3932_ (.A0(_1827_),
    .A1(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[35] ),
    .S(_1849_),
    .X(_1853_));
 sky130_fd_sc_hd__clkbuf_1 _3933_ (.A(_1853_),
    .X(_0350_));
 sky130_fd_sc_hd__mux2_1 _3934_ (.A0(_1829_),
    .A1(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[36] ),
    .S(_1849_),
    .X(_1854_));
 sky130_fd_sc_hd__clkbuf_1 _3935_ (.A(_1854_),
    .X(_0351_));
 sky130_fd_sc_hd__mux2_1 _3936_ (.A0(_1831_),
    .A1(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[37] ),
    .S(_1849_),
    .X(_1855_));
 sky130_fd_sc_hd__clkbuf_1 _3937_ (.A(_1855_),
    .X(_0352_));
 sky130_fd_sc_hd__mux2_1 _3938_ (.A0(_1833_),
    .A1(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[38] ),
    .S(_1849_),
    .X(_1856_));
 sky130_fd_sc_hd__clkbuf_1 _3939_ (.A(_1856_),
    .X(_0353_));
 sky130_fd_sc_hd__mux2_1 _3940_ (.A0(_1835_),
    .A1(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[39] ),
    .S(_1849_),
    .X(_1857_));
 sky130_fd_sc_hd__clkbuf_1 _3941_ (.A(_1857_),
    .X(_0354_));
 sky130_fd_sc_hd__nor2_1 _3942_ (.A(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_last_q[3] ),
    .B(_1807_),
    .Y(_1858_));
 sky130_fd_sc_hd__and3_1 _3943_ (.A(_1665_),
    .B(_1818_),
    .C(_1858_),
    .X(_1859_));
 sky130_fd_sc_hd__clkbuf_4 _3944_ (.A(_1859_),
    .X(_1860_));
 sky130_fd_sc_hd__mux2_1 _3945_ (.A0(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[40] ),
    .A1(\usb2uart.u_uart.uart_rx_inst.m_axis_tdata_reg[0] ),
    .S(_1860_),
    .X(_1861_));
 sky130_fd_sc_hd__clkbuf_1 _3946_ (.A(_1861_),
    .X(_0355_));
 sky130_fd_sc_hd__mux2_1 _3947_ (.A0(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[41] ),
    .A1(\usb2uart.u_uart.uart_rx_inst.m_axis_tdata_reg[1] ),
    .S(_1860_),
    .X(_1862_));
 sky130_fd_sc_hd__clkbuf_1 _3948_ (.A(_1862_),
    .X(_0356_));
 sky130_fd_sc_hd__mux2_1 _3949_ (.A0(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[42] ),
    .A1(\usb2uart.u_uart.uart_rx_inst.m_axis_tdata_reg[2] ),
    .S(_1860_),
    .X(_1863_));
 sky130_fd_sc_hd__clkbuf_1 _3950_ (.A(_1863_),
    .X(_0357_));
 sky130_fd_sc_hd__mux2_1 _3951_ (.A0(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[43] ),
    .A1(\usb2uart.u_uart.uart_rx_inst.m_axis_tdata_reg[3] ),
    .S(_1860_),
    .X(_1864_));
 sky130_fd_sc_hd__clkbuf_1 _3952_ (.A(_1864_),
    .X(_0358_));
 sky130_fd_sc_hd__mux2_1 _3953_ (.A0(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[44] ),
    .A1(\usb2uart.u_uart.uart_rx_inst.m_axis_tdata_reg[4] ),
    .S(_1860_),
    .X(_1865_));
 sky130_fd_sc_hd__clkbuf_1 _3954_ (.A(_1865_),
    .X(_0359_));
 sky130_fd_sc_hd__mux2_1 _3955_ (.A0(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[45] ),
    .A1(\usb2uart.u_uart.uart_rx_inst.m_axis_tdata_reg[5] ),
    .S(_1860_),
    .X(_1866_));
 sky130_fd_sc_hd__clkbuf_1 _3956_ (.A(_1866_),
    .X(_0360_));
 sky130_fd_sc_hd__mux2_1 _3957_ (.A0(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[46] ),
    .A1(\usb2uart.u_uart.uart_rx_inst.m_axis_tdata_reg[6] ),
    .S(_1860_),
    .X(_1867_));
 sky130_fd_sc_hd__clkbuf_1 _3958_ (.A(_1867_),
    .X(_0361_));
 sky130_fd_sc_hd__mux2_1 _3959_ (.A0(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[47] ),
    .A1(\usb2uart.u_uart.uart_rx_inst.m_axis_tdata_reg[7] ),
    .S(_1860_),
    .X(_1868_));
 sky130_fd_sc_hd__clkbuf_1 _3960_ (.A(_1868_),
    .X(_0362_));
 sky130_fd_sc_hd__nand2_1 _3961_ (.A(_1665_),
    .B(_1858_),
    .Y(_1869_));
 sky130_fd_sc_hd__or2_1 _3962_ (.A(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_last_q[0] ),
    .B(_1869_),
    .X(_1870_));
 sky130_fd_sc_hd__clkbuf_4 _3963_ (.A(_1870_),
    .X(_1871_));
 sky130_fd_sc_hd__mux2_1 _3964_ (.A0(_1819_),
    .A1(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[48] ),
    .S(_1871_),
    .X(_1872_));
 sky130_fd_sc_hd__clkbuf_1 _3965_ (.A(_1872_),
    .X(_0363_));
 sky130_fd_sc_hd__mux2_1 _3966_ (.A0(_1823_),
    .A1(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[49] ),
    .S(_1871_),
    .X(_1873_));
 sky130_fd_sc_hd__clkbuf_1 _3967_ (.A(_1873_),
    .X(_0364_));
 sky130_fd_sc_hd__mux2_1 _3968_ (.A0(_1825_),
    .A1(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[50] ),
    .S(_1871_),
    .X(_1874_));
 sky130_fd_sc_hd__clkbuf_1 _3969_ (.A(_1874_),
    .X(_0365_));
 sky130_fd_sc_hd__mux2_1 _3970_ (.A0(_1827_),
    .A1(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[51] ),
    .S(_1871_),
    .X(_1875_));
 sky130_fd_sc_hd__clkbuf_1 _3971_ (.A(_1875_),
    .X(_0366_));
 sky130_fd_sc_hd__mux2_1 _3972_ (.A0(_1829_),
    .A1(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[52] ),
    .S(_1871_),
    .X(_1876_));
 sky130_fd_sc_hd__clkbuf_1 _3973_ (.A(_1876_),
    .X(_0367_));
 sky130_fd_sc_hd__mux2_1 _3974_ (.A0(_1831_),
    .A1(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[53] ),
    .S(_1871_),
    .X(_1877_));
 sky130_fd_sc_hd__clkbuf_1 _3975_ (.A(_1877_),
    .X(_0368_));
 sky130_fd_sc_hd__mux2_1 _3976_ (.A0(_1833_),
    .A1(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[54] ),
    .S(_1871_),
    .X(_1878_));
 sky130_fd_sc_hd__clkbuf_1 _3977_ (.A(_1878_),
    .X(_0369_));
 sky130_fd_sc_hd__mux2_1 _3978_ (.A0(_1835_),
    .A1(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[55] ),
    .S(_1871_),
    .X(_1879_));
 sky130_fd_sc_hd__clkbuf_1 _3979_ (.A(_1879_),
    .X(_0370_));
 sky130_fd_sc_hd__nand3_2 _3980_ (.A(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_last_q[3] ),
    .B(_1665_),
    .C(_1805_),
    .Y(_1880_));
 sky130_fd_sc_hd__a22oi_4 _3981_ (.A1(_1804_),
    .A2(_1837_),
    .B1(_1869_),
    .B2(_1880_),
    .Y(_1881_));
 sky130_fd_sc_hd__a21o_1 _3982_ (.A1(_1869_),
    .A2(_1880_),
    .B1(_1837_),
    .X(_1882_));
 sky130_fd_sc_hd__buf_2 _3983_ (.A(_1882_),
    .X(_1883_));
 sky130_fd_sc_hd__a32o_1 _3984_ (.A1(\usb2uart.u_uart.uart_rx_inst.m_axis_tdata_reg[0] ),
    .A2(_1810_),
    .A3(_1881_),
    .B1(_1883_),
    .B2(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[56] ),
    .X(_0371_));
 sky130_fd_sc_hd__a32o_1 _3985_ (.A1(\usb2uart.u_uart.uart_rx_inst.m_axis_tdata_reg[1] ),
    .A2(_1810_),
    .A3(_1881_),
    .B1(_1883_),
    .B2(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[57] ),
    .X(_0372_));
 sky130_fd_sc_hd__a32o_1 _3986_ (.A1(\usb2uart.u_uart.uart_rx_inst.m_axis_tdata_reg[2] ),
    .A2(_1810_),
    .A3(_1881_),
    .B1(_1883_),
    .B2(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[58] ),
    .X(_0373_));
 sky130_fd_sc_hd__a32o_1 _3987_ (.A1(\usb2uart.u_uart.uart_rx_inst.m_axis_tdata_reg[3] ),
    .A2(_1810_),
    .A3(_1881_),
    .B1(_1883_),
    .B2(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[59] ),
    .X(_0374_));
 sky130_fd_sc_hd__a32o_1 _3988_ (.A1(\usb2uart.u_uart.uart_rx_inst.m_axis_tdata_reg[4] ),
    .A2(_1810_),
    .A3(_1881_),
    .B1(_1883_),
    .B2(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[60] ),
    .X(_0375_));
 sky130_fd_sc_hd__a32o_1 _3989_ (.A1(\usb2uart.u_uart.uart_rx_inst.m_axis_tdata_reg[5] ),
    .A2(_1810_),
    .A3(_1881_),
    .B1(_1883_),
    .B2(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[61] ),
    .X(_0376_));
 sky130_fd_sc_hd__a32o_1 _3990_ (.A1(\usb2uart.u_uart.uart_rx_inst.m_axis_tdata_reg[6] ),
    .A2(_1810_),
    .A3(_1881_),
    .B1(_1883_),
    .B2(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[62] ),
    .X(_0377_));
 sky130_fd_sc_hd__mux2_1 _3991_ (.A0(\usb2uart.u_uart.uart_rx_inst.m_axis_tdata_reg[7] ),
    .A1(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[63] ),
    .S(_1883_),
    .X(_1884_));
 sky130_fd_sc_hd__clkbuf_1 _3992_ (.A(_1884_),
    .X(_0378_));
 sky130_fd_sc_hd__clkbuf_4 _3993_ (.A(_1880_),
    .X(_1885_));
 sky130_fd_sc_hd__a32o_1 _3994_ (.A1(_1666_),
    .A2(_1806_),
    .A3(_1819_),
    .B1(_1885_),
    .B2(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[64] ),
    .X(_0379_));
 sky130_fd_sc_hd__a32o_1 _3995_ (.A1(_1666_),
    .A2(_1806_),
    .A3(_1823_),
    .B1(_1885_),
    .B2(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[65] ),
    .X(_0380_));
 sky130_fd_sc_hd__a32o_1 _3996_ (.A1(_1666_),
    .A2(_1806_),
    .A3(_1825_),
    .B1(_1885_),
    .B2(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[66] ),
    .X(_0381_));
 sky130_fd_sc_hd__a32o_1 _3997_ (.A1(_1666_),
    .A2(_1806_),
    .A3(_1827_),
    .B1(_1885_),
    .B2(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[67] ),
    .X(_0382_));
 sky130_fd_sc_hd__a32o_1 _3998_ (.A1(_1666_),
    .A2(_1806_),
    .A3(_1829_),
    .B1(_1885_),
    .B2(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[68] ),
    .X(_0383_));
 sky130_fd_sc_hd__a32o_1 _3999_ (.A1(_1666_),
    .A2(_1806_),
    .A3(_1831_),
    .B1(_1885_),
    .B2(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[69] ),
    .X(_0384_));
 sky130_fd_sc_hd__a32o_1 _4000_ (.A1(_1666_),
    .A2(_1806_),
    .A3(_1833_),
    .B1(_1885_),
    .B2(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[70] ),
    .X(_0385_));
 sky130_fd_sc_hd__a32o_1 _4001_ (.A1(_1666_),
    .A2(_1806_),
    .A3(_1835_),
    .B1(_1885_),
    .B2(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[71] ),
    .X(_0386_));
 sky130_fd_sc_hd__o211a_1 _4002_ (.A1(_1810_),
    .A2(_1666_),
    .B1(_1801_),
    .C1(_1885_),
    .X(_0387_));
 sky130_fd_sc_hd__and3_1 _4003_ (.A(_1582_),
    .B(_1589_),
    .C(_1665_),
    .X(_1886_));
 sky130_fd_sc_hd__a21oi_1 _4004_ (.A1(_1810_),
    .A2(_1665_),
    .B1(_1589_),
    .Y(_1887_));
 sky130_fd_sc_hd__nor2_1 _4005_ (.A(_1886_),
    .B(_1887_),
    .Y(_0388_));
 sky130_fd_sc_hd__xor2_1 _4006_ (.A(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_last_q[2] ),
    .B(_1886_),
    .X(_0389_));
 sky130_fd_sc_hd__a21bo_1 _4007_ (.A1(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_last_q[2] ),
    .A2(_1886_),
    .B1_N(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_last_q[3] ),
    .X(_1888_));
 sky130_fd_sc_hd__a21boi_1 _4008_ (.A1(_1883_),
    .A2(_1888_),
    .B1_N(_1885_),
    .Y(_0390_));
 sky130_fd_sc_hd__nor2_1 _4009_ (.A(_0951_),
    .B(_1701_),
    .Y(_0391_));
 sky130_fd_sc_hd__inv_2 _4010_ (.A(\usb2uart.u_uart.uart_tx_inst.prescale_reg[1] ),
    .Y(_1889_));
 sky130_fd_sc_hd__a21oi_1 _4011_ (.A1(_1889_),
    .A2(_1701_),
    .B1(net4),
    .Y(_1890_));
 sky130_fd_sc_hd__o21a_1 _4012_ (.A1(_1889_),
    .A2(_1701_),
    .B1(_1890_),
    .X(_0392_));
 sky130_fd_sc_hd__clkbuf_4 _4013_ (.A(_0950_),
    .X(_1891_));
 sky130_fd_sc_hd__or3_1 _4014_ (.A(\usb2uart.u_uart.uart_tx_inst.prescale_reg[2] ),
    .B(\usb2uart.u_uart.uart_tx_inst.prescale_reg[1] ),
    .C(\usb2uart.u_uart.uart_tx_inst.prescale_reg[0] ),
    .X(_1892_));
 sky130_fd_sc_hd__o21ai_1 _4015_ (.A1(\usb2uart.u_uart.uart_tx_inst.prescale_reg[1] ),
    .A2(\usb2uart.u_uart.uart_tx_inst.prescale_reg[0] ),
    .B1(\usb2uart.u_uart.uart_tx_inst.prescale_reg[2] ),
    .Y(_1893_));
 sky130_fd_sc_hd__a21o_1 _4016_ (.A1(_1892_),
    .A2(_1893_),
    .B1(_1694_),
    .X(_1894_));
 sky130_fd_sc_hd__nand2_1 _4017_ (.A(_1699_),
    .B(_1894_),
    .Y(_1895_));
 sky130_fd_sc_hd__and3_1 _4018_ (.A(_1891_),
    .B(_1698_),
    .C(_1895_),
    .X(_1896_));
 sky130_fd_sc_hd__clkbuf_1 _4019_ (.A(_1896_),
    .X(_0393_));
 sky130_fd_sc_hd__nand2_1 _4020_ (.A(\usb2uart.u_uart.uart_tx_inst.prescale_reg[3] ),
    .B(_1892_),
    .Y(_1897_));
 sky130_fd_sc_hd__nand2_1 _4021_ (.A(_1687_),
    .B(_1897_),
    .Y(_1898_));
 sky130_fd_sc_hd__and3_1 _4022_ (.A(_1891_),
    .B(_1699_),
    .C(_1898_),
    .X(_1899_));
 sky130_fd_sc_hd__clkbuf_1 _4023_ (.A(_1899_),
    .X(_0394_));
 sky130_fd_sc_hd__or2_1 _4024_ (.A(\usb2uart.u_uart.uart_tx_inst.prescale_reg[4] ),
    .B(_1687_),
    .X(_1900_));
 sky130_fd_sc_hd__nand2_1 _4025_ (.A(\usb2uart.u_uart.uart_tx_inst.prescale_reg[4] ),
    .B(_1687_),
    .Y(_1901_));
 sky130_fd_sc_hd__or2_1 _4026_ (.A(net4),
    .B(_1694_),
    .X(_1902_));
 sky130_fd_sc_hd__buf_2 _4027_ (.A(_1902_),
    .X(_1903_));
 sky130_fd_sc_hd__a21oi_1 _4028_ (.A1(_1900_),
    .A2(_1901_),
    .B1(_1903_),
    .Y(_0395_));
 sky130_fd_sc_hd__nor2_1 _4029_ (.A(\usb2uart.u_uart.uart_tx_inst.prescale_reg[4] ),
    .B(_1687_),
    .Y(_1904_));
 sky130_fd_sc_hd__a21oi_1 _4030_ (.A1(_1904_),
    .A2(_1698_),
    .B1(\usb2uart.u_uart.uart_tx_inst.prescale_reg[5] ),
    .Y(_1905_));
 sky130_fd_sc_hd__a31o_1 _4031_ (.A1(\usb2uart.u_uart.uart_tx_inst.prescale_reg[5] ),
    .A2(_1904_),
    .A3(_1698_),
    .B1(net4),
    .X(_1906_));
 sky130_fd_sc_hd__nor2_1 _4032_ (.A(_1905_),
    .B(_1906_),
    .Y(_0396_));
 sky130_fd_sc_hd__o21ai_1 _4033_ (.A1(\usb2uart.u_uart.uart_tx_inst.prescale_reg[5] ),
    .A2(_1900_),
    .B1(\usb2uart.u_uart.uart_tx_inst.prescale_reg[6] ),
    .Y(_1907_));
 sky130_fd_sc_hd__a21oi_1 _4034_ (.A1(_1688_),
    .A2(_1907_),
    .B1(_1903_),
    .Y(_0397_));
 sky130_fd_sc_hd__and2b_1 _4035_ (.A_N(_1688_),
    .B(_1698_),
    .X(_1908_));
 sky130_fd_sc_hd__xnor2_1 _4036_ (.A(\usb2uart.u_uart.uart_tx_inst.prescale_reg[7] ),
    .B(_1908_),
    .Y(_1909_));
 sky130_fd_sc_hd__nor2_1 _4037_ (.A(_0951_),
    .B(_1909_),
    .Y(_0398_));
 sky130_fd_sc_hd__or3b_1 _4038_ (.A(\usb2uart.u_uart.uart_tx_inst.prescale_reg[7] ),
    .B(_1688_),
    .C_N(_1698_),
    .X(_1910_));
 sky130_fd_sc_hd__xor2_1 _4039_ (.A(\usb2uart.u_uart.uart_tx_inst.prescale_reg[8] ),
    .B(_1910_),
    .X(_1911_));
 sky130_fd_sc_hd__nor2_1 _4040_ (.A(_0951_),
    .B(_1911_),
    .Y(_0399_));
 sky130_fd_sc_hd__or3_1 _4041_ (.A(\usb2uart.u_uart.uart_tx_inst.prescale_reg[9] ),
    .B(_1688_),
    .C(_1689_),
    .X(_1912_));
 sky130_fd_sc_hd__o21ai_1 _4042_ (.A1(_1688_),
    .A2(_1689_),
    .B1(\usb2uart.u_uart.uart_tx_inst.prescale_reg[9] ),
    .Y(_1913_));
 sky130_fd_sc_hd__a21oi_1 _4043_ (.A1(_1912_),
    .A2(_1913_),
    .B1(_1903_),
    .Y(_0400_));
 sky130_fd_sc_hd__nand2_1 _4044_ (.A(\usb2uart.u_uart.uart_tx_inst.prescale_reg[10] ),
    .B(_1912_),
    .Y(_1914_));
 sky130_fd_sc_hd__a21oi_1 _4045_ (.A1(_1690_),
    .A2(_1914_),
    .B1(_1903_),
    .Y(_0401_));
 sky130_fd_sc_hd__nor2_1 _4046_ (.A(\usb2uart.u_uart.uart_tx_inst.prescale_reg[11] ),
    .B(_1690_),
    .Y(_1915_));
 sky130_fd_sc_hd__and2_1 _4047_ (.A(\usb2uart.u_uart.uart_tx_inst.prescale_reg[11] ),
    .B(_1690_),
    .X(_1916_));
 sky130_fd_sc_hd__o211a_1 _4048_ (.A1(_1915_),
    .A2(_1916_),
    .B1(_1697_),
    .C1(_0044_),
    .X(_0402_));
 sky130_fd_sc_hd__xnor2_1 _4049_ (.A(\usb2uart.u_uart.uart_tx_inst.prescale_reg[12] ),
    .B(_1915_),
    .Y(_1917_));
 sky130_fd_sc_hd__nor2_1 _4050_ (.A(_1903_),
    .B(_1917_),
    .Y(_0403_));
 sky130_fd_sc_hd__o31ai_1 _4051_ (.A1(\usb2uart.u_uart.uart_tx_inst.prescale_reg[12] ),
    .A2(\usb2uart.u_uart.uart_tx_inst.prescale_reg[11] ),
    .A3(_1690_),
    .B1(\usb2uart.u_uart.uart_tx_inst.prescale_reg[13] ),
    .Y(_1918_));
 sky130_fd_sc_hd__a21oi_1 _4052_ (.A1(_1691_),
    .A2(_1918_),
    .B1(_1903_),
    .Y(_0404_));
 sky130_fd_sc_hd__nor2_1 _4053_ (.A(\usb2uart.u_uart.uart_tx_inst.prescale_reg[14] ),
    .B(_1691_),
    .Y(_1919_));
 sky130_fd_sc_hd__and2_1 _4054_ (.A(\usb2uart.u_uart.uart_tx_inst.prescale_reg[14] ),
    .B(_1691_),
    .X(_1920_));
 sky130_fd_sc_hd__o211a_1 _4055_ (.A1(_1919_),
    .A2(_1920_),
    .B1(_1697_),
    .C1(_0044_),
    .X(_0405_));
 sky130_fd_sc_hd__xnor2_1 _4056_ (.A(\usb2uart.u_uart.uart_tx_inst.prescale_reg[15] ),
    .B(_1919_),
    .Y(_1921_));
 sky130_fd_sc_hd__nor2_1 _4057_ (.A(_1903_),
    .B(_1921_),
    .Y(_0406_));
 sky130_fd_sc_hd__o31ai_1 _4058_ (.A1(\usb2uart.u_uart.uart_tx_inst.prescale_reg[15] ),
    .A2(\usb2uart.u_uart.uart_tx_inst.prescale_reg[14] ),
    .A3(_1691_),
    .B1(\usb2uart.u_uart.uart_tx_inst.prescale_reg[16] ),
    .Y(_1922_));
 sky130_fd_sc_hd__a21oi_1 _4059_ (.A1(_1692_),
    .A2(_1922_),
    .B1(_1903_),
    .Y(_0407_));
 sky130_fd_sc_hd__nand2_1 _4060_ (.A(\usb2uart.u_uart.uart_tx_inst.prescale_reg[17] ),
    .B(_1692_),
    .Y(_1923_));
 sky130_fd_sc_hd__a21oi_1 _4061_ (.A1(_1693_),
    .A2(_1923_),
    .B1(_1903_),
    .Y(_0408_));
 sky130_fd_sc_hd__and3_1 _4062_ (.A(\usb2uart.u_uart.uart_tx_inst.prescale_reg[18] ),
    .B(_1891_),
    .C(_1693_),
    .X(_1924_));
 sky130_fd_sc_hd__clkbuf_1 _4063_ (.A(_1924_),
    .X(_0409_));
 sky130_fd_sc_hd__or2_1 _4064_ (.A(\usb2uart.u_uart.uart_tx_inst.bit_cnt[0] ),
    .B(_1696_),
    .X(_1925_));
 sky130_fd_sc_hd__o22ai_1 _4065_ (.A1(_1682_),
    .A2(_1903_),
    .B1(_1925_),
    .B2(_0951_),
    .Y(_0410_));
 sky130_fd_sc_hd__nand2_1 _4066_ (.A(\usb2uart.u_uart.uart_tx_inst.bit_cnt[1] ),
    .B(_1925_),
    .Y(_1926_));
 sky130_fd_sc_hd__or2_1 _4067_ (.A(\usb2uart.u_uart.uart_tx_inst.bit_cnt[1] ),
    .B(_1925_),
    .X(_1927_));
 sky130_fd_sc_hd__a211oi_1 _4068_ (.A1(_1926_),
    .A2(_1927_),
    .B1(net4),
    .C1(_1683_),
    .Y(_0411_));
 sky130_fd_sc_hd__nand2_1 _4069_ (.A(\usb2uart.u_uart.uart_tx_inst.bit_cnt[2] ),
    .B(_1927_),
    .Y(_1928_));
 sky130_fd_sc_hd__or3b_1 _4070_ (.A(\usb2uart.u_uart.uart_tx_inst.bit_cnt[2] ),
    .B(_1927_),
    .C_N(\usb2uart.u_uart.uart_tx_inst.bit_cnt[3] ),
    .X(_1929_));
 sky130_fd_sc_hd__a21oi_1 _4071_ (.A1(_1928_),
    .A2(_1929_),
    .B1(_0951_),
    .Y(_0412_));
 sky130_fd_sc_hd__o21bai_1 _4072_ (.A1(\usb2uart.u_uart.uart_tx_inst.bit_cnt[2] ),
    .A2(_1927_),
    .B1_N(\usb2uart.u_uart.uart_tx_inst.bit_cnt[3] ),
    .Y(_1930_));
 sky130_fd_sc_hd__and3_1 _4073_ (.A(_1891_),
    .B(_1929_),
    .C(_1930_),
    .X(_1931_));
 sky130_fd_sc_hd__clkbuf_1 _4074_ (.A(_1931_),
    .X(_0413_));
 sky130_fd_sc_hd__nand2_1 _4075_ (.A(_1580_),
    .B(_1669_),
    .Y(_1932_));
 sky130_fd_sc_hd__o2111a_1 _4076_ (.A1(\usb2uart.u_uart.uart_tx_inst.s_axis_tready_reg ),
    .A2(_1669_),
    .B1(_1932_),
    .C1(_1891_),
    .D1(_1694_),
    .X(_0414_));
 sky130_fd_sc_hd__o211a_1 _4077_ (.A1(\usb2uart.u_uart.uart_tx_inst.data_reg[0] ),
    .A2(_1683_),
    .B1(_1684_),
    .C1(_1694_),
    .X(_1933_));
 sky130_fd_sc_hd__a211o_1 _4078_ (.A1(net10),
    .A2(_1696_),
    .B1(_1933_),
    .C1(_0951_),
    .X(_0415_));
 sky130_fd_sc_hd__or2b_1 _4079_ (.A(_1663_),
    .B_N(\usb2uart.u_uart.uart_rx_inst.m_axis_tvalid_reg ),
    .X(_1934_));
 sky130_fd_sc_hd__nand3b_4 _4080_ (.A_N(_1098_),
    .B(_1091_),
    .C(\usb2uart.u_uart.uart_rx_inst.rxd_reg ),
    .Y(_1935_));
 sky130_fd_sc_hd__a21oi_1 _4081_ (.A1(_1934_),
    .A2(_1935_),
    .B1(_0951_),
    .Y(_0416_));
 sky130_fd_sc_hd__or3_1 _4082_ (.A(_2081_),
    .B(_0498_),
    .C(_0736_),
    .X(_1936_));
 sky130_fd_sc_hd__o21ai_1 _4083_ (.A1(\usb2uart.u_usb_cdc.u_ctrl_endp.req_q[7] ),
    .A2(\usb2uart.u_usb_cdc.u_ctrl_endp.in_endp_q ),
    .B1(_0516_),
    .Y(_1937_));
 sky130_fd_sc_hd__o41a_1 _4084_ (.A1(_2017_),
    .A2(_0646_),
    .A3(_1936_),
    .A4(_1937_),
    .B1(\usb2uart.u_usb_cdc.u_sie.datain_toggle_q[1] ),
    .X(_1938_));
 sky130_fd_sc_hd__clkinv_2 _4085_ (.A(_0979_),
    .Y(_1939_));
 sky130_fd_sc_hd__nor2_1 _4086_ (.A(_0589_),
    .B(_0861_),
    .Y(_1940_));
 sky130_fd_sc_hd__and4_1 _4087_ (.A(_0588_),
    .B(_0516_),
    .C(_1940_),
    .D(_1058_),
    .X(_1941_));
 sky130_fd_sc_hd__mux2_1 _4088_ (.A0(_1938_),
    .A1(_1939_),
    .S(_1941_),
    .X(_1942_));
 sky130_fd_sc_hd__clkbuf_1 _4089_ (.A(_1942_),
    .X(_0417_));
 sky130_fd_sc_hd__and3b_1 _4090_ (.A_N(_1098_),
    .B(_1091_),
    .C(\usb2uart.u_uart.uart_rx_inst.rxd_reg ),
    .X(_1943_));
 sky130_fd_sc_hd__or2_1 _4091_ (.A(\usb2uart.u_uart.uart_rx_inst.m_axis_tdata_reg[0] ),
    .B(_1943_),
    .X(_1944_));
 sky130_fd_sc_hd__o211a_1 _4092_ (.A1(\usb2uart.u_uart.uart_rx_inst.data_reg[0] ),
    .A2(_1935_),
    .B1(_1944_),
    .C1(_0044_),
    .X(_0418_));
 sky130_fd_sc_hd__or2_1 _4093_ (.A(\usb2uart.u_uart.uart_rx_inst.m_axis_tdata_reg[1] ),
    .B(_1943_),
    .X(_1945_));
 sky130_fd_sc_hd__o211a_1 _4094_ (.A1(\usb2uart.u_uart.uart_rx_inst.data_reg[1] ),
    .A2(_1935_),
    .B1(_1945_),
    .C1(_0044_),
    .X(_0419_));
 sky130_fd_sc_hd__or2_1 _4095_ (.A(\usb2uart.u_uart.uart_rx_inst.m_axis_tdata_reg[2] ),
    .B(_1943_),
    .X(_1946_));
 sky130_fd_sc_hd__o211a_1 _4096_ (.A1(\usb2uart.u_uart.uart_rx_inst.data_reg[2] ),
    .A2(_1935_),
    .B1(_1946_),
    .C1(_0044_),
    .X(_0420_));
 sky130_fd_sc_hd__or2_1 _4097_ (.A(\usb2uart.u_uart.uart_rx_inst.m_axis_tdata_reg[3] ),
    .B(_1943_),
    .X(_1947_));
 sky130_fd_sc_hd__o211a_1 _4098_ (.A1(\usb2uart.u_uart.uart_rx_inst.data_reg[3] ),
    .A2(_1935_),
    .B1(_1947_),
    .C1(_0044_),
    .X(_0421_));
 sky130_fd_sc_hd__or2_1 _4099_ (.A(\usb2uart.u_uart.uart_rx_inst.m_axis_tdata_reg[4] ),
    .B(_1943_),
    .X(_1948_));
 sky130_fd_sc_hd__o211a_1 _4100_ (.A1(\usb2uart.u_uart.uart_rx_inst.data_reg[4] ),
    .A2(_1935_),
    .B1(_1948_),
    .C1(_0044_),
    .X(_0422_));
 sky130_fd_sc_hd__or2_1 _4101_ (.A(\usb2uart.u_uart.uart_rx_inst.m_axis_tdata_reg[5] ),
    .B(_1943_),
    .X(_1949_));
 sky130_fd_sc_hd__o211a_1 _4102_ (.A1(\usb2uart.u_uart.uart_rx_inst.data_reg[5] ),
    .A2(_1935_),
    .B1(_1949_),
    .C1(_0044_),
    .X(_0423_));
 sky130_fd_sc_hd__or2_1 _4103_ (.A(\usb2uart.u_uart.uart_rx_inst.m_axis_tdata_reg[6] ),
    .B(_1943_),
    .X(_1950_));
 sky130_fd_sc_hd__o211a_1 _4104_ (.A1(\usb2uart.u_uart.uart_rx_inst.data_reg[6] ),
    .A2(_1935_),
    .B1(_1950_),
    .C1(_0044_),
    .X(_0424_));
 sky130_fd_sc_hd__or2_1 _4105_ (.A(\usb2uart.u_uart.uart_rx_inst.m_axis_tdata_reg[7] ),
    .B(_1943_),
    .X(_1951_));
 sky130_fd_sc_hd__o211a_1 _4106_ (.A1(\usb2uart.u_uart.uart_rx_inst.data_reg[7] ),
    .A2(_1935_),
    .B1(_1951_),
    .C1(_1891_),
    .X(_0425_));
 sky130_fd_sc_hd__or2_1 _4107_ (.A(net4),
    .B(net3),
    .X(_1952_));
 sky130_fd_sc_hd__clkbuf_1 _4108_ (.A(_1952_),
    .X(_0426_));
 sky130_fd_sc_hd__nor2_2 _4109_ (.A(\usb2uart.u_uart.uart_rx_inst.prescale_reg[18] ),
    .B(_1088_),
    .Y(_1953_));
 sky130_fd_sc_hd__and2_1 _4110_ (.A(\usb2uart.u_uart.uart_rx_inst.rxd_reg ),
    .B(_1094_),
    .X(_1954_));
 sky130_fd_sc_hd__or3_2 _4111_ (.A(_1100_),
    .B(_1090_),
    .C(_1954_),
    .X(_1955_));
 sky130_fd_sc_hd__o21a_1 _4112_ (.A1(\usb2uart.u_uart.uart_rx_inst.prescale_reg[0] ),
    .A2(_1953_),
    .B1(_1955_),
    .X(_1956_));
 sky130_fd_sc_hd__nor2_1 _4113_ (.A(_1093_),
    .B(_1956_),
    .Y(_0427_));
 sky130_fd_sc_hd__xnor2_1 _4114_ (.A(\usb2uart.u_uart.uart_rx_inst.prescale_reg[1] ),
    .B(\usb2uart.u_uart.uart_rx_inst.prescale_reg[0] ),
    .Y(_1957_));
 sky130_fd_sc_hd__nor2_1 _4115_ (.A(_1090_),
    .B(_1954_),
    .Y(_1958_));
 sky130_fd_sc_hd__a21oi_1 _4116_ (.A1(_1090_),
    .A2(_1957_),
    .B1(_1958_),
    .Y(_1959_));
 sky130_fd_sc_hd__nor2_1 _4117_ (.A(_1093_),
    .B(_1959_),
    .Y(_0428_));
 sky130_fd_sc_hd__or3_1 _4118_ (.A(\usb2uart.u_uart.uart_rx_inst.prescale_reg[2] ),
    .B(\usb2uart.u_uart.uart_rx_inst.prescale_reg[1] ),
    .C(\usb2uart.u_uart.uart_rx_inst.prescale_reg[0] ),
    .X(_1960_));
 sky130_fd_sc_hd__o21ai_1 _4119_ (.A1(\usb2uart.u_uart.uart_rx_inst.prescale_reg[1] ),
    .A2(\usb2uart.u_uart.uart_rx_inst.prescale_reg[0] ),
    .B1(\usb2uart.u_uart.uart_rx_inst.prescale_reg[2] ),
    .Y(_1961_));
 sky130_fd_sc_hd__a21o_1 _4120_ (.A1(_1960_),
    .A2(_1961_),
    .B1(_1953_),
    .X(_1962_));
 sky130_fd_sc_hd__a21oi_1 _4121_ (.A1(_1955_),
    .A2(_1962_),
    .B1(_1093_),
    .Y(_0429_));
 sky130_fd_sc_hd__nand2_1 _4122_ (.A(\usb2uart.u_uart.uart_rx_inst.prescale_reg[3] ),
    .B(_1960_),
    .Y(_1963_));
 sky130_fd_sc_hd__nand2_4 _4123_ (.A(_0950_),
    .B(_1090_),
    .Y(_1964_));
 sky130_fd_sc_hd__a21oi_1 _4124_ (.A1(_1083_),
    .A2(_1963_),
    .B1(_1964_),
    .Y(_0430_));
 sky130_fd_sc_hd__xor2_1 _4125_ (.A(\usb2uart.u_uart.uart_rx_inst.prescale_reg[4] ),
    .B(_1083_),
    .X(_1965_));
 sky130_fd_sc_hd__nand2_1 _4126_ (.A(_1100_),
    .B(_1953_),
    .Y(_1966_));
 sky130_fd_sc_hd__o21a_1 _4127_ (.A1(_1953_),
    .A2(_1965_),
    .B1(_1966_),
    .X(_1967_));
 sky130_fd_sc_hd__nor2_1 _4128_ (.A(_1093_),
    .B(_1967_),
    .Y(_0431_));
 sky130_fd_sc_hd__or3_1 _4129_ (.A(\usb2uart.u_uart.uart_rx_inst.prescale_reg[5] ),
    .B(\usb2uart.u_uart.uart_rx_inst.prescale_reg[4] ),
    .C(_1083_),
    .X(_1968_));
 sky130_fd_sc_hd__o21ai_1 _4130_ (.A1(\usb2uart.u_uart.uart_rx_inst.prescale_reg[4] ),
    .A2(_1083_),
    .B1(\usb2uart.u_uart.uart_rx_inst.prescale_reg[5] ),
    .Y(_1969_));
 sky130_fd_sc_hd__a21o_1 _4131_ (.A1(_1968_),
    .A2(_1969_),
    .B1(_1953_),
    .X(_1970_));
 sky130_fd_sc_hd__a21oi_1 _4132_ (.A1(_1955_),
    .A2(_1970_),
    .B1(_1093_),
    .Y(_0432_));
 sky130_fd_sc_hd__nand2_1 _4133_ (.A(\usb2uart.u_uart.uart_rx_inst.prescale_reg[6] ),
    .B(_1968_),
    .Y(_1971_));
 sky130_fd_sc_hd__a21o_1 _4134_ (.A1(_1084_),
    .A2(_1971_),
    .B1(_1953_),
    .X(_1972_));
 sky130_fd_sc_hd__a21oi_1 _4135_ (.A1(_1966_),
    .A2(_1972_),
    .B1(_1093_),
    .Y(_0433_));
 sky130_fd_sc_hd__xnor2_1 _4136_ (.A(\usb2uart.u_uart.uart_rx_inst.prescale_reg[7] ),
    .B(_1084_),
    .Y(_1973_));
 sky130_fd_sc_hd__a21oi_1 _4137_ (.A1(_1090_),
    .A2(_1973_),
    .B1(_1958_),
    .Y(_1974_));
 sky130_fd_sc_hd__nor2_1 _4138_ (.A(_1093_),
    .B(_1974_),
    .Y(_0434_));
 sky130_fd_sc_hd__or3_1 _4139_ (.A(\usb2uart.u_uart.uart_rx_inst.prescale_reg[8] ),
    .B(\usb2uart.u_uart.uart_rx_inst.prescale_reg[7] ),
    .C(_1084_),
    .X(_1975_));
 sky130_fd_sc_hd__o21ai_1 _4140_ (.A1(\usb2uart.u_uart.uart_rx_inst.prescale_reg[7] ),
    .A2(_1084_),
    .B1(\usb2uart.u_uart.uart_rx_inst.prescale_reg[8] ),
    .Y(_1976_));
 sky130_fd_sc_hd__a21o_1 _4141_ (.A1(_1975_),
    .A2(_1976_),
    .B1(_1953_),
    .X(_1977_));
 sky130_fd_sc_hd__a21oi_1 _4142_ (.A1(_1955_),
    .A2(_1977_),
    .B1(_1093_),
    .Y(_0435_));
 sky130_fd_sc_hd__nand2_1 _4143_ (.A(\usb2uart.u_uart.uart_rx_inst.prescale_reg[9] ),
    .B(_1975_),
    .Y(_1978_));
 sky130_fd_sc_hd__a21oi_1 _4144_ (.A1(_1085_),
    .A2(_1978_),
    .B1(_1964_),
    .Y(_0436_));
 sky130_fd_sc_hd__nor2_1 _4145_ (.A(\usb2uart.u_uart.uart_rx_inst.prescale_reg[10] ),
    .B(_1085_),
    .Y(_1979_));
 sky130_fd_sc_hd__and2_1 _4146_ (.A(\usb2uart.u_uart.uart_rx_inst.prescale_reg[10] ),
    .B(_1085_),
    .X(_1980_));
 sky130_fd_sc_hd__o211a_1 _4147_ (.A1(_1979_),
    .A2(_1980_),
    .B1(_1090_),
    .C1(_1891_),
    .X(_0437_));
 sky130_fd_sc_hd__xnor2_1 _4148_ (.A(\usb2uart.u_uart.uart_rx_inst.prescale_reg[11] ),
    .B(_1979_),
    .Y(_1981_));
 sky130_fd_sc_hd__nor2_1 _4149_ (.A(_1964_),
    .B(_1981_),
    .Y(_0438_));
 sky130_fd_sc_hd__o31ai_1 _4150_ (.A1(\usb2uart.u_uart.uart_rx_inst.prescale_reg[11] ),
    .A2(\usb2uart.u_uart.uart_rx_inst.prescale_reg[10] ),
    .A3(_1085_),
    .B1(\usb2uart.u_uart.uart_rx_inst.prescale_reg[12] ),
    .Y(_1982_));
 sky130_fd_sc_hd__a21oi_1 _4151_ (.A1(_1086_),
    .A2(_1982_),
    .B1(_1964_),
    .Y(_0439_));
 sky130_fd_sc_hd__nor2_1 _4152_ (.A(\usb2uart.u_uart.uart_rx_inst.prescale_reg[13] ),
    .B(_1086_),
    .Y(_1983_));
 sky130_fd_sc_hd__and2_1 _4153_ (.A(\usb2uart.u_uart.uart_rx_inst.prescale_reg[13] ),
    .B(_1086_),
    .X(_1984_));
 sky130_fd_sc_hd__o211a_1 _4154_ (.A1(_1983_),
    .A2(_1984_),
    .B1(_1090_),
    .C1(_1891_),
    .X(_0440_));
 sky130_fd_sc_hd__xnor2_1 _4155_ (.A(\usb2uart.u_uart.uart_rx_inst.prescale_reg[14] ),
    .B(_1983_),
    .Y(_1985_));
 sky130_fd_sc_hd__nor2_1 _4156_ (.A(_1964_),
    .B(_1985_),
    .Y(_0441_));
 sky130_fd_sc_hd__o31ai_1 _4157_ (.A1(\usb2uart.u_uart.uart_rx_inst.prescale_reg[14] ),
    .A2(\usb2uart.u_uart.uart_rx_inst.prescale_reg[13] ),
    .A3(_1086_),
    .B1(\usb2uart.u_uart.uart_rx_inst.prescale_reg[15] ),
    .Y(_1986_));
 sky130_fd_sc_hd__a21oi_1 _4158_ (.A1(_1087_),
    .A2(_1986_),
    .B1(_1964_),
    .Y(_0442_));
 sky130_fd_sc_hd__or2_1 _4159_ (.A(\usb2uart.u_uart.uart_rx_inst.prescale_reg[16] ),
    .B(_1087_),
    .X(_1987_));
 sky130_fd_sc_hd__nand2_1 _4160_ (.A(\usb2uart.u_uart.uart_rx_inst.prescale_reg[16] ),
    .B(_1087_),
    .Y(_1988_));
 sky130_fd_sc_hd__a21oi_1 _4161_ (.A1(_1987_),
    .A2(_1988_),
    .B1(_1964_),
    .Y(_0443_));
 sky130_fd_sc_hd__o21ai_1 _4162_ (.A1(\usb2uart.u_uart.uart_rx_inst.prescale_reg[16] ),
    .A2(_1087_),
    .B1(\usb2uart.u_uart.uart_rx_inst.prescale_reg[17] ),
    .Y(_1989_));
 sky130_fd_sc_hd__a21oi_1 _4163_ (.A1(_1088_),
    .A2(_1989_),
    .B1(_1964_),
    .Y(_0444_));
 sky130_fd_sc_hd__and3_1 _4164_ (.A(\usb2uart.u_uart.uart_rx_inst.prescale_reg[18] ),
    .B(_0950_),
    .C(_1088_),
    .X(_1990_));
 sky130_fd_sc_hd__clkbuf_1 _4165_ (.A(_1990_),
    .X(_0445_));
 sky130_fd_sc_hd__mux2_1 _4166_ (.A0(_1955_),
    .A1(_1953_),
    .S(\usb2uart.u_uart.uart_rx_inst.bit_cnt[0] ),
    .X(_1991_));
 sky130_fd_sc_hd__nor2_1 _4167_ (.A(_0951_),
    .B(_1991_),
    .Y(_0446_));
 sky130_fd_sc_hd__a21oi_2 _4168_ (.A1(\usb2uart.u_uart.uart_rx_inst.rxd_reg ),
    .A2(_1100_),
    .B1(_1090_),
    .Y(_1992_));
 sky130_fd_sc_hd__and2_1 _4169_ (.A(\usb2uart.u_uart.uart_rx_inst.bit_cnt[1] ),
    .B(\usb2uart.u_uart.uart_rx_inst.bit_cnt[0] ),
    .X(_1993_));
 sky130_fd_sc_hd__nor2_1 _4170_ (.A(_1098_),
    .B(_1993_),
    .Y(_1994_));
 sky130_fd_sc_hd__o21ai_1 _4171_ (.A1(_1954_),
    .A2(_1994_),
    .B1(_1992_),
    .Y(_1995_));
 sky130_fd_sc_hd__o211a_1 _4172_ (.A1(\usb2uart.u_uart.uart_rx_inst.bit_cnt[1] ),
    .A2(_1992_),
    .B1(_1995_),
    .C1(_1891_),
    .X(_0447_));
 sky130_fd_sc_hd__xnor2_1 _4173_ (.A(\usb2uart.u_uart.uart_rx_inst.bit_cnt[2] ),
    .B(_1098_),
    .Y(_1996_));
 sky130_fd_sc_hd__o31ai_1 _4174_ (.A1(_1100_),
    .A2(_1954_),
    .A3(_1996_),
    .B1(_1992_),
    .Y(_1997_));
 sky130_fd_sc_hd__o211a_1 _4175_ (.A1(\usb2uart.u_uart.uart_rx_inst.bit_cnt[2] ),
    .A2(_1992_),
    .B1(_1997_),
    .C1(_1891_),
    .X(_0448_));
 sky130_fd_sc_hd__a21oi_1 _4176_ (.A1(_1097_),
    .A2(_1098_),
    .B1(_1954_),
    .Y(_1998_));
 sky130_fd_sc_hd__o21ai_1 _4177_ (.A1(_1090_),
    .A2(_1998_),
    .B1(\usb2uart.u_uart.uart_rx_inst.bit_cnt[3] ),
    .Y(_1999_));
 sky130_fd_sc_hd__nand2_1 _4178_ (.A(_1100_),
    .B(_1992_),
    .Y(_2000_));
 sky130_fd_sc_hd__a21oi_1 _4179_ (.A1(_1999_),
    .A2(_2000_),
    .B1(_0951_),
    .Y(_0449_));
 sky130_fd_sc_hd__dfstp_1 _4180_ (.CLK(clknet_leaf_11_user_clock2),
    .D(_0017_),
    .SET_B(net31),
    .Q(\usb2uart.u_usb_cdc.u_sie.phy_state_q[0] ));
 sky130_fd_sc_hd__dfrtp_1 _4181_ (.CLK(clknet_leaf_14_user_clock2),
    .D(_0020_),
    .RESET_B(net39),
    .Q(\usb2uart.u_usb_cdc.u_sie.phy_state_q[1] ));
 sky130_fd_sc_hd__dfrtp_1 _4182_ (.CLK(clknet_leaf_11_user_clock2),
    .D(_0021_),
    .RESET_B(net31),
    .Q(\usb2uart.u_usb_cdc.u_sie.phy_state_q[2] ));
 sky130_fd_sc_hd__dfrtp_1 _4183_ (.CLK(clknet_leaf_12_user_clock2),
    .D(_0022_),
    .RESET_B(net28),
    .Q(\usb2uart.u_usb_cdc.u_sie.phy_state_q[3] ));
 sky130_fd_sc_hd__dfrtp_2 _4184_ (.CLK(clknet_leaf_21_user_clock2),
    .D(_0023_),
    .RESET_B(net41),
    .Q(\usb2uart.u_usb_cdc.u_sie.phy_state_q[4] ));
 sky130_fd_sc_hd__dfrtp_1 _4185_ (.CLK(clknet_leaf_11_user_clock2),
    .D(_0024_),
    .RESET_B(net32),
    .Q(\usb2uart.u_usb_cdc.u_sie.phy_state_q[5] ));
 sky130_fd_sc_hd__dfrtp_1 _4186_ (.CLK(clknet_leaf_11_user_clock2),
    .D(_0025_),
    .RESET_B(net31),
    .Q(\usb2uart.u_usb_cdc.u_sie.phy_state_q[6] ));
 sky130_fd_sc_hd__dfrtp_4 _4187_ (.CLK(clknet_leaf_21_user_clock2),
    .D(_0026_),
    .RESET_B(net41),
    .Q(\usb2uart.u_usb_cdc.u_sie.phy_state_q[7] ));
 sky130_fd_sc_hd__dfrtp_1 _4188_ (.CLK(clknet_leaf_15_user_clock2),
    .D(_0027_),
    .RESET_B(net39),
    .Q(\usb2uart.u_usb_cdc.u_sie.phy_state_q[8] ));
 sky130_fd_sc_hd__dfrtp_4 _4189_ (.CLK(clknet_leaf_11_user_clock2),
    .D(_0028_),
    .RESET_B(net29),
    .Q(\usb2uart.u_usb_cdc.u_sie.phy_state_q[9] ));
 sky130_fd_sc_hd__dfrtp_2 _4190_ (.CLK(clknet_leaf_14_user_clock2),
    .D(_0018_),
    .RESET_B(net41),
    .Q(\usb2uart.u_usb_cdc.u_sie.phy_state_q[10] ));
 sky130_fd_sc_hd__dfrtp_2 _4191_ (.CLK(clknet_leaf_14_user_clock2),
    .D(_0019_),
    .RESET_B(net41),
    .Q(\usb2uart.u_usb_cdc.u_sie.phy_state_q[11] ));
 sky130_fd_sc_hd__dfstp_1 _4192_ (.CLK(clknet_leaf_13_user_clock2),
    .D(_0013_),
    .SET_B(net31),
    .Q(\usb2uart.u_usb_cdc.u_ctrl_endp.state_q[0] ));
 sky130_fd_sc_hd__dfrtp_1 _4193_ (.CLK(clknet_leaf_13_user_clock2),
    .D(_0014_),
    .RESET_B(net31),
    .Q(\usb2uart.u_usb_cdc.u_ctrl_endp.state_q[1] ));
 sky130_fd_sc_hd__dfrtp_1 _4194_ (.CLK(clknet_leaf_13_user_clock2),
    .D(_0015_),
    .RESET_B(net39),
    .Q(\usb2uart.u_usb_cdc.ctrl_stall ));
 sky130_fd_sc_hd__dfrtp_4 _4195_ (.CLK(clknet_leaf_13_user_clock2),
    .D(_0016_),
    .RESET_B(net31),
    .Q(\usb2uart.u_usb_cdc.u_ctrl_endp.state_q[3] ));
 sky130_fd_sc_hd__dfstp_4 _4196_ (.CLK(clknet_leaf_16_user_clock2),
    .D(_0034_),
    .SET_B(net43),
    .Q(net6));
 sky130_fd_sc_hd__dfrtp_2 _4197_ (.CLK(clknet_leaf_17_user_clock2),
    .D(_0035_),
    .RESET_B(net40),
    .Q(\usb2uart.u_usb_cdc.u_sie.u_phy_tx.tx_state_q[1] ));
 sky130_fd_sc_hd__dfrtp_1 _4198_ (.CLK(clknet_leaf_16_user_clock2),
    .D(_0036_),
    .RESET_B(net40),
    .Q(\usb2uart.u_usb_cdc.u_sie.u_phy_tx.tx_state_q[2] ));
 sky130_fd_sc_hd__dfrtp_4 _4199_ (.CLK(clknet_leaf_17_user_clock2),
    .D(_0037_),
    .RESET_B(net40),
    .Q(\usb2uart.u_usb_cdc.u_sie.u_phy_tx.tx_state_q[3] ));
 sky130_fd_sc_hd__dfstp_1 _4200_ (.CLK(clknet_leaf_16_user_clock2),
    .D(_0029_),
    .SET_B(net61),
    .Q(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.rx_state_q[0] ));
 sky130_fd_sc_hd__dfrtp_4 _4201_ (.CLK(clknet_leaf_15_user_clock2),
    .D(_0030_),
    .RESET_B(net60),
    .Q(\usb2uart.u_usb_cdc.u_sie.rx_err ));
 sky130_fd_sc_hd__dfrtp_2 _4202_ (.CLK(clknet_leaf_11_user_clock2),
    .D(_0031_),
    .RESET_B(net59),
    .Q(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.rx_state_q[2] ));
 sky130_fd_sc_hd__dfrtp_2 _4203_ (.CLK(clknet_leaf_10_user_clock2),
    .D(_0032_),
    .RESET_B(net59),
    .Q(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.rx_state_q[3] ));
 sky130_fd_sc_hd__dfrtp_1 _4204_ (.CLK(clknet_leaf_15_user_clock2),
    .D(_0033_),
    .RESET_B(net60),
    .Q(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.rx_state_q[4] ));
 sky130_fd_sc_hd__dfrtp_1 _4205_ (.CLK(clknet_leaf_12_user_clock2),
    .D(_0046_),
    .RESET_B(net29),
    .Q(\usb2uart.u_usb_cdc.u_sie.datain_toggle_q[0] ));
 sky130_fd_sc_hd__dfrtp_1 _4206_ (.CLK(clknet_leaf_32_user_clock2),
    .D(_0000_),
    .RESET_B(net33),
    .Q(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_state_q[1] ));
 sky130_fd_sc_hd__dfrtp_1 _4207_ (.CLK(clknet_leaf_10_user_clock2),
    .D(_0047_),
    .RESET_B(net57),
    .Q(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.cnt_q[0] ));
 sky130_fd_sc_hd__dfrtp_1 _4208_ (.CLK(clknet_leaf_9_user_clock2),
    .D(_0048_),
    .RESET_B(net55),
    .Q(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.cnt_q[1] ));
 sky130_fd_sc_hd__dfrtp_1 _4209_ (.CLK(clknet_leaf_9_user_clock2),
    .D(_0049_),
    .RESET_B(net56),
    .Q(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.cnt_q[3] ));
 sky130_fd_sc_hd__dfrtp_1 _4210_ (.CLK(clknet_leaf_9_user_clock2),
    .D(_0050_),
    .RESET_B(net56),
    .Q(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.cnt_q[4] ));
 sky130_fd_sc_hd__dfrtp_1 _4211_ (.CLK(clknet_leaf_8_user_clock2),
    .D(_0051_),
    .RESET_B(net56),
    .Q(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.cnt_q[6] ));
 sky130_fd_sc_hd__dfrtp_1 _4212_ (.CLK(clknet_leaf_8_user_clock2),
    .D(_0052_),
    .RESET_B(net55),
    .Q(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.cnt_q[7] ));
 sky130_fd_sc_hd__dfrtp_1 _4213_ (.CLK(clknet_leaf_9_user_clock2),
    .D(_0053_),
    .RESET_B(net55),
    .Q(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.cnt_q[8] ));
 sky130_fd_sc_hd__dfrtp_1 _4214_ (.CLK(clknet_leaf_8_user_clock2),
    .D(_0054_),
    .RESET_B(net55),
    .Q(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.cnt_q[9] ));
 sky130_fd_sc_hd__dfrtp_1 _4215_ (.CLK(clknet_leaf_8_user_clock2),
    .D(_0055_),
    .RESET_B(net55),
    .Q(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.cnt_q[10] ));
 sky130_fd_sc_hd__dfrtp_1 _4216_ (.CLK(clknet_leaf_8_user_clock2),
    .D(_0056_),
    .RESET_B(net55),
    .Q(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.cnt_q[11] ));
 sky130_fd_sc_hd__dfrtp_1 _4217_ (.CLK(clknet_leaf_9_user_clock2),
    .D(_0057_),
    .RESET_B(net55),
    .Q(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.cnt_q[12] ));
 sky130_fd_sc_hd__dfrtp_1 _4218_ (.CLK(clknet_leaf_10_user_clock2),
    .D(_0058_),
    .RESET_B(net55),
    .Q(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.cnt_q[13] ));
 sky130_fd_sc_hd__dfrtp_1 _4219_ (.CLK(clknet_leaf_10_user_clock2),
    .D(_0059_),
    .RESET_B(net57),
    .Q(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.cnt_q[14] ));
 sky130_fd_sc_hd__dfrtp_1 _4220_ (.CLK(clknet_leaf_9_user_clock2),
    .D(_0060_),
    .RESET_B(net55),
    .Q(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.cnt_q[15] ));
 sky130_fd_sc_hd__dfrtp_1 _4221_ (.CLK(clknet_leaf_10_user_clock2),
    .D(_0061_),
    .RESET_B(net57),
    .Q(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.cnt_q[16] ));
 sky130_fd_sc_hd__dfrtp_1 _4222_ (.CLK(clknet_leaf_10_user_clock2),
    .D(_0062_),
    .RESET_B(net57),
    .Q(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.cnt_q[17] ));
 sky130_fd_sc_hd__dfstp_1 _4223_ (.CLK(clknet_leaf_3_user_clock2),
    .D(_0001_),
    .SET_B(net24),
    .Q(\usb2uart.u_usb_cdc.u_ctrl_endp.req_q[0] ));
 sky130_fd_sc_hd__dfrtp_1 _4224_ (.CLK(clknet_leaf_4_user_clock2),
    .D(_0004_),
    .RESET_B(net21),
    .Q(\usb2uart.u_usb_cdc.u_ctrl_endp.req_q[1] ));
 sky130_fd_sc_hd__dfrtp_1 _4225_ (.CLK(clknet_leaf_3_user_clock2),
    .D(_0005_),
    .RESET_B(net27),
    .Q(\usb2uart.u_usb_cdc.u_ctrl_endp.req_q[2] ));
 sky130_fd_sc_hd__dfrtp_4 _4226_ (.CLK(clknet_leaf_4_user_clock2),
    .D(_0006_),
    .RESET_B(net21),
    .Q(\usb2uart.u_usb_cdc.u_ctrl_endp.req_q[3] ));
 sky130_fd_sc_hd__dfrtp_1 _4227_ (.CLK(clknet_leaf_2_user_clock2),
    .D(_0007_),
    .RESET_B(net24),
    .Q(\usb2uart.u_usb_cdc.u_ctrl_endp.req_q[4] ));
 sky130_fd_sc_hd__dfrtp_1 _4228_ (.CLK(clknet_leaf_4_user_clock2),
    .D(_0008_),
    .RESET_B(net17),
    .Q(\usb2uart.u_usb_cdc.u_ctrl_endp.req_q[5] ));
 sky130_fd_sc_hd__dfrtp_1 _4229_ (.CLK(clknet_leaf_4_user_clock2),
    .D(_0009_),
    .RESET_B(net28),
    .Q(\usb2uart.u_usb_cdc.u_ctrl_endp.req_q[6] ));
 sky130_fd_sc_hd__dfrtp_4 _4230_ (.CLK(clknet_leaf_4_user_clock2),
    .D(_0010_),
    .RESET_B(net28),
    .Q(\usb2uart.u_usb_cdc.u_ctrl_endp.req_q[7] ));
 sky130_fd_sc_hd__dfrtp_1 _4231_ (.CLK(clknet_leaf_3_user_clock2),
    .D(_0011_),
    .RESET_B(net27),
    .Q(\usb2uart.u_usb_cdc.u_ctrl_endp.req_q[8] ));
 sky130_fd_sc_hd__dfrtp_1 _4232_ (.CLK(clknet_leaf_5_user_clock2),
    .D(_0012_),
    .RESET_B(net17),
    .Q(\usb2uart.u_usb_cdc.u_ctrl_endp.req_q[9] ));
 sky130_fd_sc_hd__dfrtp_2 _4233_ (.CLK(clknet_leaf_3_user_clock2),
    .D(_0002_),
    .RESET_B(net25),
    .Q(\usb2uart.u_usb_cdc.u_ctrl_endp.req_q[10] ));
 sky130_fd_sc_hd__dfrtp_1 _4234_ (.CLK(clknet_leaf_1_user_clock2),
    .D(_0003_),
    .RESET_B(net17),
    .Q(\usb2uart.u_usb_cdc.u_ctrl_endp.req_q[11] ));
 sky130_fd_sc_hd__dfrtp_1 _4235_ (.CLK(clknet_leaf_16_user_clock2),
    .D(_0063_),
    .RESET_B(net40),
    .Q(\usb2uart.u_usb_cdc.u_sie.u_phy_tx.tx_valid_q ));
 sky130_fd_sc_hd__dfrtp_1 _4236_ (.CLK(clknet_leaf_30_user_clock2),
    .D(net301),
    .RESET_B(_0044_),
    .Q(\usb2uart.u_usb_cdc.rstn ));
 sky130_fd_sc_hd__dfrtp_1 _4237_ (.CLK(clknet_leaf_30_user_clock2),
    .D(net263),
    .RESET_B(_0045_),
    .Q(\usb2uart.u_usb_cdc.rstn_sq[1] ));
 sky130_fd_sc_hd__dfrtp_2 _4238_ (.CLK(clknet_leaf_17_user_clock2),
    .D(_0064_),
    .RESET_B(net50),
    .Q(\usb2uart.u_usb_cdc.u_sie.u_phy_tx.data_q[0] ));
 sky130_fd_sc_hd__dfrtp_1 _4239_ (.CLK(clknet_leaf_17_user_clock2),
    .D(_0065_),
    .RESET_B(net50),
    .Q(\usb2uart.u_usb_cdc.u_sie.u_phy_tx.data_q[1] ));
 sky130_fd_sc_hd__dfrtp_1 _4240_ (.CLK(clknet_leaf_17_user_clock2),
    .D(_0066_),
    .RESET_B(net42),
    .Q(\usb2uart.u_usb_cdc.u_sie.u_phy_tx.data_q[2] ));
 sky130_fd_sc_hd__dfrtp_1 _4241_ (.CLK(clknet_leaf_18_user_clock2),
    .D(_0067_),
    .RESET_B(net50),
    .Q(\usb2uart.u_usb_cdc.u_sie.u_phy_tx.data_q[3] ));
 sky130_fd_sc_hd__dfrtp_1 _4242_ (.CLK(clknet_leaf_18_user_clock2),
    .D(_0068_),
    .RESET_B(net51),
    .Q(\usb2uart.u_usb_cdc.u_sie.u_phy_tx.data_q[4] ));
 sky130_fd_sc_hd__dfrtp_1 _4243_ (.CLK(clknet_leaf_18_user_clock2),
    .D(_0069_),
    .RESET_B(net50),
    .Q(\usb2uart.u_usb_cdc.u_sie.u_phy_tx.data_q[5] ));
 sky130_fd_sc_hd__dfrtp_1 _4244_ (.CLK(clknet_leaf_15_user_clock2),
    .D(_0070_),
    .RESET_B(net40),
    .Q(\usb2uart.u_usb_cdc.u_sie.u_phy_tx.data_q[6] ));
 sky130_fd_sc_hd__dfstp_1 _4245_ (.CLK(clknet_leaf_17_user_clock2),
    .D(_0071_),
    .SET_B(net40),
    .Q(\usb2uart.u_usb_cdc.u_sie.u_phy_tx.data_q[7] ));
 sky130_fd_sc_hd__dfstp_1 _4246_ (.CLK(clknet_leaf_18_user_clock2),
    .D(_0072_),
    .SET_B(net52),
    .Q(\usb2uart.u_usb_cdc.u_sie.u_phy_tx.bit_cnt_q[0] ));
 sky130_fd_sc_hd__dfstp_1 _4247_ (.CLK(clknet_leaf_18_user_clock2),
    .D(_0073_),
    .SET_B(net50),
    .Q(\usb2uart.u_usb_cdc.u_sie.u_phy_tx.bit_cnt_q[1] ));
 sky130_fd_sc_hd__dfstp_1 _4248_ (.CLK(clknet_leaf_18_user_clock2),
    .D(_0074_),
    .SET_B(net50),
    .Q(\usb2uart.u_usb_cdc.u_sie.u_phy_tx.bit_cnt_q[2] ));
 sky130_fd_sc_hd__dfstp_1 _4249_ (.CLK(clknet_leaf_16_user_clock2),
    .D(_0075_),
    .SET_B(net43),
    .Q(\usb2uart.u_usb_cdc.u_sie.u_phy_tx.nrzi_q ));
 sky130_fd_sc_hd__dfrtp_1 _4250_ (.CLK(clknet_leaf_17_user_clock2),
    .D(_0076_),
    .RESET_B(net50),
    .Q(\usb2uart.u_usb_cdc.u_sie.u_phy_tx.stuffing_cnt_q[0] ));
 sky130_fd_sc_hd__dfrtp_1 _4251_ (.CLK(clknet_leaf_17_user_clock2),
    .D(_0077_),
    .RESET_B(net40),
    .Q(\usb2uart.u_usb_cdc.u_sie.u_phy_tx.stuffing_cnt_q[1] ));
 sky130_fd_sc_hd__dfrtp_1 _4252_ (.CLK(clknet_leaf_16_user_clock2),
    .D(_0078_),
    .RESET_B(net42),
    .Q(\usb2uart.u_usb_cdc.u_sie.u_phy_tx.stuffing_cnt_q[2] ));
 sky130_fd_sc_hd__dfrtp_1 _4253_ (.CLK(clknet_leaf_16_user_clock2),
    .D(_0042_),
    .RESET_B(net40),
    .Q(\usb2uart.u_usb_cdc.u_sie.u_phy_tx.clk_cnt_q[0] ));
 sky130_fd_sc_hd__dfrtp_1 _4254_ (.CLK(clknet_leaf_17_user_clock2),
    .D(_0043_),
    .RESET_B(net40),
    .Q(\usb2uart.u_usb_cdc.u_sie.u_phy_tx.clk_cnt_q[1] ));
 sky130_fd_sc_hd__dfrtp_4 _4255_ (.CLK(clknet_leaf_9_user_clock2),
    .D(_0079_),
    .RESET_B(net55),
    .Q(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.rx_en_q ));
 sky130_fd_sc_hd__dfrtp_1 _4256_ (.CLK(clknet_leaf_10_user_clock2),
    .D(_0040_),
    .RESET_B(net61),
    .Q(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.clk_cnt_q[0] ));
 sky130_fd_sc_hd__dfrtp_1 _4257_ (.CLK(clknet_leaf_10_user_clock2),
    .D(_0041_),
    .RESET_B(net58),
    .Q(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.clk_cnt_q[1] ));
 sky130_fd_sc_hd__dfrtp_1 _4258_ (.CLK(clknet_leaf_16_user_clock2),
    .D(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.dp_q[1] ),
    .RESET_B(net61),
    .Q(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.dp_q[0] ));
 sky130_fd_sc_hd__dfrtp_1 _4259_ (.CLK(clknet_leaf_16_user_clock2),
    .D(net299),
    .RESET_B(net59),
    .Q(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.dp_q[1] ));
 sky130_fd_sc_hd__dfrtp_1 _4260_ (.CLK(clknet_leaf_10_user_clock2),
    .D(net2),
    .RESET_B(net59),
    .Q(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.dp_q[2] ));
 sky130_fd_sc_hd__dfrtp_2 _4261_ (.CLK(clknet_leaf_10_user_clock2),
    .D(_0080_),
    .RESET_B(net57),
    .Q(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.cnt_q[2] ));
 sky130_fd_sc_hd__dfrtp_1 _4262_ (.CLK(clknet_leaf_9_user_clock2),
    .D(_0081_),
    .RESET_B(net57),
    .Q(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.cnt_q[5] ));
 sky130_fd_sc_hd__dfrtp_4 _4263_ (.CLK(clknet_leaf_11_user_clock2),
    .D(_0082_),
    .RESET_B(net57),
    .Q(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.rx_valid_fq ));
 sky130_fd_sc_hd__dfrtp_4 _4264_ (.CLK(clknet_leaf_11_user_clock2),
    .D(_0083_),
    .RESET_B(net59),
    .Q(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.rx_valid_fd ));
 sky130_fd_sc_hd__dfrtp_1 _4265_ (.CLK(clknet_leaf_10_user_clock2),
    .D(_0084_),
    .RESET_B(net58),
    .Q(net7));
 sky130_fd_sc_hd__dfrtp_1 _4266_ (.CLK(clknet_leaf_10_user_clock2),
    .D(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.dn_q[1] ),
    .RESET_B(net59),
    .Q(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.dn_q[0] ));
 sky130_fd_sc_hd__dfrtp_1 _4267_ (.CLK(clknet_leaf_10_user_clock2),
    .D(net300),
    .RESET_B(net59),
    .Q(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.dn_q[1] ));
 sky130_fd_sc_hd__dfrtp_1 _4268_ (.CLK(clknet_leaf_10_user_clock2),
    .D(net1),
    .RESET_B(net61),
    .Q(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.dn_q[2] ));
 sky130_fd_sc_hd__dfrtp_1 _4269_ (.CLK(clknet_leaf_13_user_clock2),
    .D(_0085_),
    .RESET_B(net39),
    .Q(\usb2uart.u_usb_cdc.u_sie.dataout_toggle_q[0] ));
 sky130_fd_sc_hd__dfrtp_4 _4270_ (.CLK(clknet_leaf_13_user_clock2),
    .D(_0086_),
    .RESET_B(net31),
    .Q(\usb2uart.u_usb_cdc.in_data_ack ));
 sky130_fd_sc_hd__dfrtp_1 _4271_ (.CLK(clknet_leaf_17_user_clock2),
    .D(_0087_),
    .RESET_B(net60),
    .Q(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.data_q[0] ));
 sky130_fd_sc_hd__dfrtp_1 _4272_ (.CLK(clknet_leaf_15_user_clock2),
    .D(_0088_),
    .RESET_B(net60),
    .Q(\usb2uart.u_usb_cdc.u_sie.rx_data[0] ));
 sky130_fd_sc_hd__dfrtp_1 _4273_ (.CLK(clknet_leaf_15_user_clock2),
    .D(_0089_),
    .RESET_B(net60),
    .Q(\usb2uart.u_usb_cdc.u_sie.rx_data[1] ));
 sky130_fd_sc_hd__dfrtp_1 _4274_ (.CLK(clknet_leaf_15_user_clock2),
    .D(_0090_),
    .RESET_B(net60),
    .Q(\usb2uart.u_usb_cdc.u_sie.rx_data[2] ));
 sky130_fd_sc_hd__dfrtp_1 _4275_ (.CLK(clknet_leaf_15_user_clock2),
    .D(_0091_),
    .RESET_B(net60),
    .Q(\usb2uart.u_usb_cdc.u_sie.rx_data[3] ));
 sky130_fd_sc_hd__dfrtp_2 _4276_ (.CLK(clknet_leaf_15_user_clock2),
    .D(_0092_),
    .RESET_B(net60),
    .Q(\usb2uart.u_usb_cdc.u_sie.rx_data[4] ));
 sky130_fd_sc_hd__dfrtp_1 _4277_ (.CLK(clknet_leaf_15_user_clock2),
    .D(_0093_),
    .RESET_B(net60),
    .Q(\usb2uart.u_usb_cdc.u_sie.rx_data[5] ));
 sky130_fd_sc_hd__dfrtp_1 _4278_ (.CLK(clknet_leaf_15_user_clock2),
    .D(_0094_),
    .RESET_B(net60),
    .Q(\usb2uart.u_usb_cdc.u_sie.rx_data[6] ));
 sky130_fd_sc_hd__dfstp_1 _4279_ (.CLK(clknet_leaf_15_user_clock2),
    .D(_0095_),
    .SET_B(net59),
    .Q(\usb2uart.u_usb_cdc.u_sie.rx_data[7] ));
 sky130_fd_sc_hd__dfrtp_1 _4280_ (.CLK(clknet_leaf_10_user_clock2),
    .D(_0096_),
    .RESET_B(net57),
    .Q(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.stuffing_cnt_q[0] ));
 sky130_fd_sc_hd__dfrtp_1 _4281_ (.CLK(clknet_leaf_11_user_clock2),
    .D(_0097_),
    .RESET_B(net57),
    .Q(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.stuffing_cnt_q[1] ));
 sky130_fd_sc_hd__dfrtp_1 _4282_ (.CLK(clknet_leaf_11_user_clock2),
    .D(_0098_),
    .RESET_B(net57),
    .Q(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.stuffing_cnt_q[2] ));
 sky130_fd_sc_hd__dfrtp_1 _4283_ (.CLK(clknet_leaf_16_user_clock2),
    .D(_0099_),
    .RESET_B(net61),
    .Q(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.nrzi_q[0] ));
 sky130_fd_sc_hd__dfrtp_1 _4284_ (.CLK(clknet_leaf_10_user_clock2),
    .D(_0100_),
    .RESET_B(net59),
    .Q(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.nrzi_q[1] ));
 sky130_fd_sc_hd__dfrtp_2 _4285_ (.CLK(clknet_leaf_16_user_clock2),
    .D(_0101_),
    .RESET_B(net61),
    .Q(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.nrzi_q[2] ));
 sky130_fd_sc_hd__dfrtp_2 _4286_ (.CLK(clknet_leaf_10_user_clock2),
    .D(_0102_),
    .RESET_B(net59),
    .Q(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.nrzi_q[3] ));
 sky130_fd_sc_hd__dfxtp_1 _4287_ (.CLK(clknet_leaf_27_user_clock2),
    .D(_0103_),
    .Q(\usb2uart.u_uart.uart_rx_inst.data_reg[0] ));
 sky130_fd_sc_hd__dfxtp_1 _4288_ (.CLK(clknet_leaf_30_user_clock2),
    .D(_0104_),
    .Q(\usb2uart.u_uart.uart_rx_inst.data_reg[1] ));
 sky130_fd_sc_hd__dfxtp_1 _4289_ (.CLK(clknet_leaf_30_user_clock2),
    .D(_0105_),
    .Q(\usb2uart.u_uart.uart_rx_inst.data_reg[2] ));
 sky130_fd_sc_hd__dfxtp_1 _4290_ (.CLK(clknet_leaf_30_user_clock2),
    .D(_0106_),
    .Q(\usb2uart.u_uart.uart_rx_inst.data_reg[3] ));
 sky130_fd_sc_hd__dfxtp_1 _4291_ (.CLK(clknet_leaf_30_user_clock2),
    .D(_0107_),
    .Q(\usb2uart.u_uart.uart_rx_inst.data_reg[4] ));
 sky130_fd_sc_hd__dfxtp_1 _4292_ (.CLK(clknet_leaf_30_user_clock2),
    .D(_0108_),
    .Q(\usb2uart.u_uart.uart_rx_inst.data_reg[5] ));
 sky130_fd_sc_hd__dfxtp_1 _4293_ (.CLK(clknet_leaf_29_user_clock2),
    .D(_0109_),
    .Q(\usb2uart.u_uart.uart_rx_inst.data_reg[6] ));
 sky130_fd_sc_hd__dfxtp_1 _4294_ (.CLK(clknet_leaf_30_user_clock2),
    .D(_0110_),
    .Q(\usb2uart.u_uart.uart_rx_inst.data_reg[7] ));
 sky130_fd_sc_hd__dfrtp_1 _4295_ (.CLK(clknet_leaf_15_user_clock2),
    .D(_0111_),
    .RESET_B(net41),
    .Q(\usb2uart.u_usb_cdc.u_sie.pid_q[0] ));
 sky130_fd_sc_hd__dfrtp_1 _4296_ (.CLK(clknet_leaf_15_user_clock2),
    .D(_0112_),
    .RESET_B(net39),
    .Q(\usb2uart.u_usb_cdc.u_sie.pid_q[1] ));
 sky130_fd_sc_hd__dfrtp_1 _4297_ (.CLK(clknet_leaf_15_user_clock2),
    .D(_0113_),
    .RESET_B(net39),
    .Q(\usb2uart.u_usb_cdc.u_sie.pid_q[2] ));
 sky130_fd_sc_hd__dfrtp_4 _4298_ (.CLK(clknet_leaf_15_user_clock2),
    .D(_0114_),
    .RESET_B(net39),
    .Q(\usb2uart.u_usb_cdc.u_sie.pid_q[3] ));
 sky130_fd_sc_hd__dfrtp_1 _4299_ (.CLK(clknet_leaf_6_user_clock2),
    .D(_0115_),
    .RESET_B(net19),
    .Q(\usb2uart.u_usb_cdc.u_sie.addr_q[0] ));
 sky130_fd_sc_hd__dfrtp_1 _4300_ (.CLK(clknet_leaf_6_user_clock2),
    .D(_0116_),
    .RESET_B(net20),
    .Q(\usb2uart.u_usb_cdc.u_sie.addr_q[1] ));
 sky130_fd_sc_hd__dfrtp_1 _4301_ (.CLK(clknet_leaf_6_user_clock2),
    .D(_0117_),
    .RESET_B(net19),
    .Q(\usb2uart.u_usb_cdc.u_sie.addr_q[2] ));
 sky130_fd_sc_hd__dfrtp_1 _4302_ (.CLK(clknet_leaf_6_user_clock2),
    .D(_0118_),
    .RESET_B(net19),
    .Q(\usb2uart.u_usb_cdc.u_sie.addr_q[3] ));
 sky130_fd_sc_hd__dfrtp_1 _4303_ (.CLK(clknet_leaf_6_user_clock2),
    .D(_0119_),
    .RESET_B(net19),
    .Q(\usb2uart.u_usb_cdc.u_sie.addr_q[4] ));
 sky130_fd_sc_hd__dfrtp_1 _4304_ (.CLK(clknet_leaf_6_user_clock2),
    .D(_0120_),
    .RESET_B(net19),
    .Q(\usb2uart.u_usb_cdc.u_sie.addr_q[5] ));
 sky130_fd_sc_hd__dfrtp_1 _4305_ (.CLK(clknet_leaf_6_user_clock2),
    .D(_0121_),
    .RESET_B(net20),
    .Q(\usb2uart.u_usb_cdc.u_sie.addr_q[6] ));
 sky130_fd_sc_hd__dfrtp_1 _4306_ (.CLK(clknet_leaf_13_user_clock2),
    .D(_0122_),
    .RESET_B(net39),
    .Q(\usb2uart.u_usb_cdc.u_sie.dataout_toggle_q[1] ));
 sky130_fd_sc_hd__dfrtp_1 _4307_ (.CLK(clknet_leaf_20_user_clock2),
    .D(_0123_),
    .RESET_B(net51),
    .Q(\usb2uart.u_usb_cdc.u_sie.in_byte_q[0] ));
 sky130_fd_sc_hd__dfrtp_1 _4308_ (.CLK(clknet_leaf_20_user_clock2),
    .D(_0124_),
    .RESET_B(net51),
    .Q(\usb2uart.u_usb_cdc.u_sie.in_byte_q[1] ));
 sky130_fd_sc_hd__dfrtp_1 _4309_ (.CLK(clknet_leaf_21_user_clock2),
    .D(_0125_),
    .RESET_B(net41),
    .Q(\usb2uart.u_usb_cdc.u_sie.in_byte_q[2] ));
 sky130_fd_sc_hd__dfrtp_1 _4310_ (.CLK(clknet_leaf_21_user_clock2),
    .D(_0126_),
    .RESET_B(net41),
    .Q(\usb2uart.u_usb_cdc.u_sie.in_byte_q[3] ));
 sky130_fd_sc_hd__dfrtp_1 _4311_ (.CLK(clknet_leaf_12_user_clock2),
    .D(_0127_),
    .RESET_B(net28),
    .Q(\usb2uart.u_usb_cdc.u_sie.delay_cnt_q[0] ));
 sky130_fd_sc_hd__dfrtp_1 _4312_ (.CLK(clknet_leaf_11_user_clock2),
    .D(_0128_),
    .RESET_B(net30),
    .Q(\usb2uart.u_usb_cdc.u_sie.delay_cnt_q[1] ));
 sky130_fd_sc_hd__dfrtp_1 _4313_ (.CLK(clknet_leaf_9_user_clock2),
    .D(_0129_),
    .RESET_B(net30),
    .Q(\usb2uart.u_usb_cdc.u_sie.delay_cnt_q[2] ));
 sky130_fd_sc_hd__dfrtp_1 _4314_ (.CLK(clknet_leaf_11_user_clock2),
    .D(_0130_),
    .RESET_B(net31),
    .Q(\usb2uart.u_usb_cdc.u_sie.delay_cnt_q[3] ));
 sky130_fd_sc_hd__dfrtp_1 _4315_ (.CLK(clknet_leaf_11_user_clock2),
    .D(_0131_),
    .RESET_B(net30),
    .Q(\usb2uart.u_usb_cdc.u_sie.delay_cnt_q[4] ));
 sky130_fd_sc_hd__dfrtp_1 _4316_ (.CLK(clknet_leaf_12_user_clock2),
    .D(_0132_),
    .RESET_B(net31),
    .Q(\usb2uart.u_usb_cdc.u_sie.out_eop_q ));
 sky130_fd_sc_hd__dfrtp_1 _4317_ (.CLK(clknet_leaf_19_user_clock2),
    .D(_0133_),
    .RESET_B(net52),
    .Q(\usb2uart.u_usb_cdc.u_sie.crc16_q[0] ));
 sky130_fd_sc_hd__dfrtp_1 _4318_ (.CLK(clknet_leaf_19_user_clock2),
    .D(_0134_),
    .RESET_B(net52),
    .Q(\usb2uart.u_usb_cdc.u_sie.crc16_q[1] ));
 sky130_fd_sc_hd__dfrtp_1 _4319_ (.CLK(clknet_leaf_19_user_clock2),
    .D(_0135_),
    .RESET_B(net52),
    .Q(\usb2uart.u_usb_cdc.u_sie.crc16_q[2] ));
 sky130_fd_sc_hd__dfrtp_1 _4320_ (.CLK(clknet_leaf_19_user_clock2),
    .D(_0136_),
    .RESET_B(net51),
    .Q(\usb2uart.u_usb_cdc.u_sie.crc16_q[3] ));
 sky130_fd_sc_hd__dfrtp_1 _4321_ (.CLK(clknet_leaf_19_user_clock2),
    .D(_0137_),
    .RESET_B(net52),
    .Q(\usb2uart.u_usb_cdc.u_sie.crc16_q[4] ));
 sky130_fd_sc_hd__dfrtp_1 _4322_ (.CLK(clknet_leaf_19_user_clock2),
    .D(_0138_),
    .RESET_B(net50),
    .Q(\usb2uart.u_usb_cdc.u_sie.crc16_q[5] ));
 sky130_fd_sc_hd__dfrtp_1 _4323_ (.CLK(clknet_leaf_18_user_clock2),
    .D(_0139_),
    .RESET_B(net52),
    .Q(\usb2uart.u_usb_cdc.u_sie.crc16_q[6] ));
 sky130_fd_sc_hd__dfrtp_1 _4324_ (.CLK(clknet_leaf_19_user_clock2),
    .D(_0140_),
    .RESET_B(net51),
    .Q(\usb2uart.u_usb_cdc.u_sie.crc16_q[7] ));
 sky130_fd_sc_hd__dfrtp_1 _4325_ (.CLK(clknet_leaf_19_user_clock2),
    .D(_0141_),
    .RESET_B(net52),
    .Q(\usb2uart.u_usb_cdc.u_sie.crc16_q[8] ));
 sky130_fd_sc_hd__dfrtp_1 _4326_ (.CLK(clknet_leaf_20_user_clock2),
    .D(_0142_),
    .RESET_B(net51),
    .Q(\usb2uart.u_usb_cdc.u_sie.crc16_q[9] ));
 sky130_fd_sc_hd__dfrtp_1 _4327_ (.CLK(clknet_leaf_15_user_clock2),
    .D(_0143_),
    .RESET_B(net42),
    .Q(\usb2uart.u_usb_cdc.u_sie.crc16_q[10] ));
 sky130_fd_sc_hd__dfrtp_1 _4328_ (.CLK(clknet_leaf_17_user_clock2),
    .D(_0144_),
    .RESET_B(net50),
    .Q(\usb2uart.u_usb_cdc.u_sie.crc16_q[11] ));
 sky130_fd_sc_hd__dfrtp_1 _4329_ (.CLK(clknet_leaf_19_user_clock2),
    .D(_0145_),
    .RESET_B(net50),
    .Q(\usb2uart.u_usb_cdc.u_sie.crc16_q[12] ));
 sky130_fd_sc_hd__dfrtp_1 _4330_ (.CLK(clknet_leaf_15_user_clock2),
    .D(_0146_),
    .RESET_B(net40),
    .Q(\usb2uart.u_usb_cdc.u_sie.crc16_q[13] ));
 sky130_fd_sc_hd__dfrtp_1 _4331_ (.CLK(clknet_leaf_17_user_clock2),
    .D(_0147_),
    .RESET_B(net42),
    .Q(\usb2uart.u_usb_cdc.u_sie.crc16_q[14] ));
 sky130_fd_sc_hd__dfrtp_1 _4332_ (.CLK(clknet_leaf_19_user_clock2),
    .D(_0148_),
    .RESET_B(net51),
    .Q(\usb2uart.u_usb_cdc.u_sie.crc16_q[15] ));
 sky130_fd_sc_hd__dfrtp_4 _4333_ (.CLK(clknet_leaf_12_user_clock2),
    .D(_0149_),
    .RESET_B(net29),
    .Q(\usb2uart.u_usb_cdc.endp[0] ));
 sky130_fd_sc_hd__dfrtp_1 _4334_ (.CLK(clknet_leaf_12_user_clock2),
    .D(_0150_),
    .RESET_B(net28),
    .Q(\usb2uart.u_usb_cdc.endp[1] ));
 sky130_fd_sc_hd__dfrtp_1 _4335_ (.CLK(clknet_leaf_12_user_clock2),
    .D(_0151_),
    .RESET_B(net28),
    .Q(\usb2uart.u_usb_cdc.endp[2] ));
 sky130_fd_sc_hd__dfrtp_1 _4336_ (.CLK(clknet_leaf_12_user_clock2),
    .D(_0152_),
    .RESET_B(net28),
    .Q(\usb2uart.u_usb_cdc.endp[3] ));
 sky130_fd_sc_hd__dfrtp_2 _4337_ (.CLK(clknet_leaf_4_user_clock2),
    .D(_0153_),
    .RESET_B(net62),
    .Q(\usb2uart.u_usb_cdc.u_ctrl_endp.dev_state_qq[0] ));
 sky130_fd_sc_hd__dfrtp_4 _4338_ (.CLK(clknet_leaf_4_user_clock2),
    .D(_0154_),
    .RESET_B(net62),
    .Q(\usb2uart.u_usb_cdc.u_ctrl_endp.dev_state_qq[1] ));
 sky130_fd_sc_hd__dfrtp_1 _4339_ (.CLK(clknet_leaf_13_user_clock2),
    .D(_0155_),
    .RESET_B(net31),
    .Q(\usb2uart.u_usb_cdc.out_err ));
 sky130_fd_sc_hd__dfrtp_1 _4340_ (.CLK(clknet_leaf_20_user_clock2),
    .D(_0156_),
    .RESET_B(net51),
    .Q(\usb2uart.u_usb_cdc.u_sie.data_q[0] ));
 sky130_fd_sc_hd__dfrtp_2 _4341_ (.CLK(clknet_leaf_14_user_clock2),
    .D(_0157_),
    .RESET_B(net41),
    .Q(\usb2uart.u_usb_cdc.u_sie.data_q[1] ));
 sky130_fd_sc_hd__dfrtp_4 _4342_ (.CLK(clknet_leaf_14_user_clock2),
    .D(_0158_),
    .RESET_B(net43),
    .Q(\usb2uart.u_usb_cdc.u_sie.data_q[2] ));
 sky130_fd_sc_hd__dfrtp_1 _4343_ (.CLK(clknet_leaf_13_user_clock2),
    .D(_0159_),
    .RESET_B(net39),
    .Q(\usb2uart.u_usb_cdc.u_sie.data_q[3] ));
 sky130_fd_sc_hd__dfrtp_4 _4344_ (.CLK(clknet_leaf_21_user_clock2),
    .D(_0160_),
    .RESET_B(net41),
    .Q(\usb2uart.u_usb_cdc.u_sie.data_q[4] ));
 sky130_fd_sc_hd__dfrtp_4 _4345_ (.CLK(clknet_leaf_20_user_clock2),
    .D(_0161_),
    .RESET_B(net41),
    .Q(\usb2uart.u_usb_cdc.u_sie.data_q[5] ));
 sky130_fd_sc_hd__dfrtp_4 _4346_ (.CLK(clknet_leaf_20_user_clock2),
    .D(_0162_),
    .RESET_B(net51),
    .Q(\usb2uart.u_usb_cdc.u_sie.data_q[6] ));
 sky130_fd_sc_hd__dfrtp_4 _4347_ (.CLK(clknet_leaf_14_user_clock2),
    .D(_0163_),
    .RESET_B(net39),
    .Q(\usb2uart.u_usb_cdc.u_sie.data_q[7] ));
 sky130_fd_sc_hd__dfrtp_2 _4348_ (.CLK(clknet_2_1__leaf_user_clock2),
    .D(_0164_),
    .RESET_B(net21),
    .Q(\usb2uart.u_usb_cdc.out_data[0] ));
 sky130_fd_sc_hd__dfrtp_4 _4349_ (.CLK(clknet_leaf_12_user_clock2),
    .D(_0165_),
    .RESET_B(net28),
    .Q(\usb2uart.u_usb_cdc.out_data[1] ));
 sky130_fd_sc_hd__dfrtp_4 _4350_ (.CLK(clknet_leaf_4_user_clock2),
    .D(_0166_),
    .RESET_B(net21),
    .Q(\usb2uart.u_usb_cdc.out_data[2] ));
 sky130_fd_sc_hd__dfrtp_4 _4351_ (.CLK(clknet_leaf_4_user_clock2),
    .D(_0167_),
    .RESET_B(net21),
    .Q(\usb2uart.u_usb_cdc.out_data[3] ));
 sky130_fd_sc_hd__dfrtp_4 _4352_ (.CLK(clknet_leaf_4_user_clock2),
    .D(_0168_),
    .RESET_B(net21),
    .Q(\usb2uart.u_usb_cdc.out_data[4] ));
 sky130_fd_sc_hd__dfrtp_4 _4353_ (.CLK(clknet_leaf_4_user_clock2),
    .D(_0169_),
    .RESET_B(net21),
    .Q(\usb2uart.u_usb_cdc.out_data[5] ));
 sky130_fd_sc_hd__dfrtp_1 _4354_ (.CLK(clknet_leaf_4_user_clock2),
    .D(_0170_),
    .RESET_B(net22),
    .Q(\usb2uart.u_usb_cdc.out_data[6] ));
 sky130_fd_sc_hd__dfrtp_4 _4355_ (.CLK(clknet_leaf_4_user_clock2),
    .D(_0171_),
    .RESET_B(net28),
    .Q(\usb2uart.u_usb_cdc.out_data[7] ));
 sky130_fd_sc_hd__dfrtp_1 _4356_ (.CLK(clknet_leaf_5_user_clock2),
    .D(_0172_),
    .RESET_B(net13),
    .Q(\usb2uart.u_usb_cdc.u_ctrl_endp.rec_q[0] ));
 sky130_fd_sc_hd__dfrtp_1 _4357_ (.CLK(clknet_leaf_5_user_clock2),
    .D(_0173_),
    .RESET_B(net13),
    .Q(\usb2uart.u_usb_cdc.u_ctrl_endp.rec_q[1] ));
 sky130_fd_sc_hd__dfrtp_1 _4358_ (.CLK(clknet_leaf_4_user_clock2),
    .D(_0174_),
    .RESET_B(net29),
    .Q(\usb2uart.u_usb_cdc.u_ctrl_endp.in_endp_q ));
 sky130_fd_sc_hd__dfstp_1 _4359_ (.CLK(clknet_leaf_4_user_clock2),
    .D(_0175_),
    .SET_B(net21),
    .Q(\usb2uart.u_usb_cdc.u_ctrl_endp.dev_state_q[0] ));
 sky130_fd_sc_hd__dfrtp_1 _4360_ (.CLK(clknet_leaf_4_user_clock2),
    .D(_0176_),
    .RESET_B(net28),
    .Q(\usb2uart.u_usb_cdc.u_ctrl_endp.dev_state_q[1] ));
 sky130_fd_sc_hd__dfrtp_4 _4361_ (.CLK(clknet_leaf_32_user_clock2),
    .D(_0177_),
    .RESET_B(net34),
    .Q(\usb2uart.u_usb_cdc.bulk_out_nak ));
 sky130_fd_sc_hd__dfrtp_1 _4362_ (.CLK(clknet_leaf_6_user_clock2),
    .D(_0178_),
    .RESET_B(net13),
    .Q(\usb2uart.u_usb_cdc.u_ctrl_endp.addr_q[0] ));
 sky130_fd_sc_hd__dfrtp_1 _4363_ (.CLK(clknet_leaf_4_user_clock2),
    .D(_0179_),
    .RESET_B(net21),
    .Q(\usb2uart.u_usb_cdc.u_ctrl_endp.addr_q[1] ));
 sky130_fd_sc_hd__dfrtp_1 _4364_ (.CLK(clknet_leaf_6_user_clock2),
    .D(_0180_),
    .RESET_B(net19),
    .Q(\usb2uart.u_usb_cdc.u_ctrl_endp.addr_q[2] ));
 sky130_fd_sc_hd__dfrtp_1 _4365_ (.CLK(clknet_leaf_5_user_clock2),
    .D(_0181_),
    .RESET_B(net20),
    .Q(\usb2uart.u_usb_cdc.u_ctrl_endp.addr_q[3] ));
 sky130_fd_sc_hd__dfrtp_1 _4366_ (.CLK(clknet_leaf_5_user_clock2),
    .D(_0182_),
    .RESET_B(net13),
    .Q(\usb2uart.u_usb_cdc.u_ctrl_endp.addr_q[4] ));
 sky130_fd_sc_hd__dfrtp_1 _4367_ (.CLK(clknet_leaf_6_user_clock2),
    .D(_0183_),
    .RESET_B(net19),
    .Q(\usb2uart.u_usb_cdc.u_ctrl_endp.addr_q[5] ));
 sky130_fd_sc_hd__dfrtp_1 _4368_ (.CLK(clknet_leaf_5_user_clock2),
    .D(_0184_),
    .RESET_B(net13),
    .Q(\usb2uart.u_usb_cdc.u_ctrl_endp.addr_q[6] ));
 sky130_fd_sc_hd__dfrtp_2 _4369_ (.CLK(clknet_leaf_32_user_clock2),
    .D(_0185_),
    .RESET_B(net34),
    .Q(\usb2uart.u_usb_cdc.u_ctrl_endp.byte_cnt_q[0] ));
 sky130_fd_sc_hd__dfrtp_4 _4370_ (.CLK(clknet_leaf_32_user_clock2),
    .D(_0186_),
    .RESET_B(net34),
    .Q(\usb2uart.u_usb_cdc.u_ctrl_endp.byte_cnt_q[1] ));
 sky130_fd_sc_hd__dfrtp_2 _4371_ (.CLK(clknet_leaf_32_user_clock2),
    .D(_0187_),
    .RESET_B(net34),
    .Q(\usb2uart.u_usb_cdc.u_ctrl_endp.byte_cnt_q[2] ));
 sky130_fd_sc_hd__dfrtp_2 _4372_ (.CLK(clknet_leaf_32_user_clock2),
    .D(_0188_),
    .RESET_B(net34),
    .Q(\usb2uart.u_usb_cdc.u_ctrl_endp.byte_cnt_q[3] ));
 sky130_fd_sc_hd__dfrtp_1 _4373_ (.CLK(clknet_leaf_22_user_clock2),
    .D(_0189_),
    .RESET_B(net34),
    .Q(\usb2uart.u_usb_cdc.u_ctrl_endp.byte_cnt_q[4] ));
 sky130_fd_sc_hd__dfrtp_2 _4374_ (.CLK(clknet_leaf_22_user_clock2),
    .D(_0190_),
    .RESET_B(net37),
    .Q(\usb2uart.u_usb_cdc.u_ctrl_endp.byte_cnt_q[5] ));
 sky130_fd_sc_hd__dfrtp_4 _4375_ (.CLK(clknet_leaf_22_user_clock2),
    .D(_0191_),
    .RESET_B(net37),
    .Q(\usb2uart.u_usb_cdc.u_ctrl_endp.byte_cnt_q[6] ));
 sky130_fd_sc_hd__dfrtp_1 _4376_ (.CLK(clknet_leaf_3_user_clock2),
    .D(_0192_),
    .RESET_B(net27),
    .Q(\usb2uart.u_usb_cdc.u_ctrl_endp.max_length_q[0] ));
 sky130_fd_sc_hd__dfrtp_1 _4377_ (.CLK(clknet_leaf_3_user_clock2),
    .D(_0193_),
    .RESET_B(net24),
    .Q(\usb2uart.u_usb_cdc.u_ctrl_endp.max_length_q[1] ));
 sky130_fd_sc_hd__dfrtp_1 _4378_ (.CLK(clknet_leaf_3_user_clock2),
    .D(_0194_),
    .RESET_B(net27),
    .Q(\usb2uart.u_usb_cdc.u_ctrl_endp.max_length_q[2] ));
 sky130_fd_sc_hd__dfrtp_1 _4379_ (.CLK(clknet_leaf_3_user_clock2),
    .D(_0195_),
    .RESET_B(net27),
    .Q(\usb2uart.u_usb_cdc.u_ctrl_endp.max_length_q[3] ));
 sky130_fd_sc_hd__dfrtp_1 _4380_ (.CLK(clknet_leaf_3_user_clock2),
    .D(_0196_),
    .RESET_B(net27),
    .Q(\usb2uart.u_usb_cdc.u_ctrl_endp.max_length_q[4] ));
 sky130_fd_sc_hd__dfrtp_1 _4381_ (.CLK(clknet_leaf_3_user_clock2),
    .D(_0197_),
    .RESET_B(net27),
    .Q(\usb2uart.u_usb_cdc.u_ctrl_endp.max_length_q[5] ));
 sky130_fd_sc_hd__dfrtp_1 _4382_ (.CLK(clknet_leaf_3_user_clock2),
    .D(_0198_),
    .RESET_B(net25),
    .Q(\usb2uart.u_usb_cdc.u_ctrl_endp.max_length_q[6] ));
 sky130_fd_sc_hd__dfrtp_2 _4383_ (.CLK(clknet_leaf_2_user_clock2),
    .D(_0199_),
    .RESET_B(net24),
    .Q(\usb2uart.u_usb_cdc.u_ctrl_endp.in_dir_q ));
 sky130_fd_sc_hd__dfrtp_2 _4384_ (.CLK(clknet_leaf_5_user_clock2),
    .D(_0200_),
    .RESET_B(net14),
    .Q(\usb2uart.u_usb_cdc.u_ctrl_endp.class_q ));
 sky130_fd_sc_hd__dfrtp_1 _4385_ (.CLK(clknet_leaf_6_user_clock2),
    .D(_0201_),
    .RESET_B(net20),
    .Q(\usb2uart.u_usb_cdc.addr[0] ));
 sky130_fd_sc_hd__dfrtp_1 _4386_ (.CLK(clknet_leaf_4_user_clock2),
    .D(_0202_),
    .RESET_B(net21),
    .Q(\usb2uart.u_usb_cdc.addr[1] ));
 sky130_fd_sc_hd__dfrtp_1 _4387_ (.CLK(clknet_leaf_6_user_clock2),
    .D(_0203_),
    .RESET_B(net19),
    .Q(\usb2uart.u_usb_cdc.addr[2] ));
 sky130_fd_sc_hd__dfrtp_1 _4388_ (.CLK(clknet_leaf_6_user_clock2),
    .D(_0204_),
    .RESET_B(net20),
    .Q(\usb2uart.u_usb_cdc.addr[3] ));
 sky130_fd_sc_hd__dfrtp_1 _4389_ (.CLK(clknet_leaf_6_user_clock2),
    .D(_0205_),
    .RESET_B(net19),
    .Q(\usb2uart.u_usb_cdc.addr[4] ));
 sky130_fd_sc_hd__dfrtp_1 _4390_ (.CLK(clknet_leaf_6_user_clock2),
    .D(_0206_),
    .RESET_B(net20),
    .Q(\usb2uart.u_usb_cdc.addr[5] ));
 sky130_fd_sc_hd__dfrtp_1 _4391_ (.CLK(clknet_leaf_6_user_clock2),
    .D(_0207_),
    .RESET_B(net19),
    .Q(\usb2uart.u_usb_cdc.addr[6] ));
 sky130_fd_sc_hd__dfrtp_1 _4392_ (.CLK(clknet_leaf_21_user_clock2),
    .D(\usb2uart.u_usb_cdc.ctrl_in_req ),
    .RESET_B(net62),
    .Q(\usb2uart.u_usb_cdc.u_ctrl_endp.in_req_q ));
 sky130_fd_sc_hd__dfrtp_4 _4393_ (.CLK(clknet_leaf_9_user_clock2),
    .D(_0039_),
    .RESET_B(net56),
    .Q(\usb2uart.u_usb_cdc.u_ctrl_endp.usb_reset_q ));
 sky130_fd_sc_hd__dfrtp_1 _4394_ (.CLK(clknet_leaf_32_user_clock2),
    .D(_0208_),
    .RESET_B(net26),
    .Q(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_last_qq[0] ));
 sky130_fd_sc_hd__dfrtp_1 _4395_ (.CLK(clknet_leaf_32_user_clock2),
    .D(_0209_),
    .RESET_B(net27),
    .Q(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_last_qq[1] ));
 sky130_fd_sc_hd__dfrtp_4 _4396_ (.CLK(clknet_leaf_32_user_clock2),
    .D(_0210_),
    .RESET_B(net34),
    .Q(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_last_qq[2] ));
 sky130_fd_sc_hd__dfrtp_1 _4397_ (.CLK(clknet_leaf_32_user_clock2),
    .D(_0211_),
    .RESET_B(net27),
    .Q(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_last_qq[3] ));
 sky130_fd_sc_hd__dfrtp_1 _4398_ (.CLK(clknet_leaf_33_user_clock2),
    .D(_0212_),
    .RESET_B(net26),
    .Q(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_last_q[0] ));
 sky130_fd_sc_hd__dfrtp_1 _4399_ (.CLK(clknet_leaf_32_user_clock2),
    .D(_0213_),
    .RESET_B(net33),
    .Q(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_last_q[1] ));
 sky130_fd_sc_hd__dfrtp_1 _4400_ (.CLK(clknet_leaf_32_user_clock2),
    .D(_0214_),
    .RESET_B(net33),
    .Q(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_last_q[2] ));
 sky130_fd_sc_hd__dfrtp_1 _4401_ (.CLK(clknet_leaf_32_user_clock2),
    .D(_0215_),
    .RESET_B(net26),
    .Q(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_last_q[3] ));
 sky130_fd_sc_hd__dfrtp_1 _4402_ (.CLK(clknet_leaf_1_user_clock2),
    .D(_0216_),
    .RESET_B(net17),
    .Q(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[0] ));
 sky130_fd_sc_hd__dfrtp_1 _4403_ (.CLK(clknet_leaf_2_user_clock2),
    .D(_0217_),
    .RESET_B(net24),
    .Q(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[1] ));
 sky130_fd_sc_hd__dfrtp_1 _4404_ (.CLK(clknet_leaf_0_user_clock2),
    .D(_0218_),
    .RESET_B(net13),
    .Q(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[2] ));
 sky130_fd_sc_hd__dfrtp_1 _4405_ (.CLK(clknet_leaf_1_user_clock2),
    .D(_0219_),
    .RESET_B(net13),
    .Q(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[3] ));
 sky130_fd_sc_hd__dfrtp_1 _4406_ (.CLK(clknet_leaf_1_user_clock2),
    .D(_0220_),
    .RESET_B(net14),
    .Q(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[4] ));
 sky130_fd_sc_hd__dfrtp_1 _4407_ (.CLK(clknet_leaf_1_user_clock2),
    .D(_0221_),
    .RESET_B(net17),
    .Q(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[5] ));
 sky130_fd_sc_hd__dfrtp_1 _4408_ (.CLK(clknet_leaf_1_user_clock2),
    .D(_0222_),
    .RESET_B(net18),
    .Q(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[6] ));
 sky130_fd_sc_hd__dfrtp_1 _4409_ (.CLK(clknet_leaf_3_user_clock2),
    .D(_0223_),
    .RESET_B(net24),
    .Q(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[7] ));
 sky130_fd_sc_hd__dfrtp_1 _4410_ (.CLK(clknet_leaf_1_user_clock2),
    .D(_0224_),
    .RESET_B(net17),
    .Q(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[8] ));
 sky130_fd_sc_hd__dfrtp_1 _4411_ (.CLK(clknet_leaf_2_user_clock2),
    .D(_0225_),
    .RESET_B(net24),
    .Q(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[9] ));
 sky130_fd_sc_hd__dfrtp_1 _4412_ (.CLK(clknet_leaf_1_user_clock2),
    .D(_0226_),
    .RESET_B(net14),
    .Q(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[10] ));
 sky130_fd_sc_hd__dfrtp_1 _4413_ (.CLK(clknet_leaf_1_user_clock2),
    .D(_0227_),
    .RESET_B(net14),
    .Q(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[11] ));
 sky130_fd_sc_hd__dfrtp_1 _4414_ (.CLK(clknet_leaf_1_user_clock2),
    .D(_0228_),
    .RESET_B(net14),
    .Q(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[12] ));
 sky130_fd_sc_hd__dfrtp_1 _4415_ (.CLK(clknet_leaf_1_user_clock2),
    .D(_0229_),
    .RESET_B(net17),
    .Q(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[13] ));
 sky130_fd_sc_hd__dfrtp_1 _4416_ (.CLK(clknet_leaf_1_user_clock2),
    .D(_0230_),
    .RESET_B(net17),
    .Q(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[14] ));
 sky130_fd_sc_hd__dfrtp_1 _4417_ (.CLK(clknet_leaf_2_user_clock2),
    .D(_0231_),
    .RESET_B(net24),
    .Q(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[15] ));
 sky130_fd_sc_hd__dfrtp_1 _4418_ (.CLK(clknet_leaf_0_user_clock2),
    .D(_0232_),
    .RESET_B(net15),
    .Q(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[16] ));
 sky130_fd_sc_hd__dfrtp_1 _4419_ (.CLK(clknet_leaf_2_user_clock2),
    .D(_0233_),
    .RESET_B(net23),
    .Q(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[17] ));
 sky130_fd_sc_hd__dfrtp_1 _4420_ (.CLK(clknet_leaf_0_user_clock2),
    .D(_0234_),
    .RESET_B(net13),
    .Q(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[18] ));
 sky130_fd_sc_hd__dfrtp_1 _4421_ (.CLK(clknet_leaf_0_user_clock2),
    .D(_0235_),
    .RESET_B(net13),
    .Q(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[19] ));
 sky130_fd_sc_hd__dfrtp_1 _4422_ (.CLK(clknet_leaf_0_user_clock2),
    .D(_0236_),
    .RESET_B(net11),
    .Q(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[20] ));
 sky130_fd_sc_hd__dfrtp_1 _4423_ (.CLK(clknet_leaf_1_user_clock2),
    .D(_0237_),
    .RESET_B(net16),
    .Q(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[21] ));
 sky130_fd_sc_hd__dfrtp_1 _4424_ (.CLK(clknet_leaf_1_user_clock2),
    .D(_0238_),
    .RESET_B(net17),
    .Q(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[22] ));
 sky130_fd_sc_hd__dfrtp_1 _4425_ (.CLK(clknet_leaf_2_user_clock2),
    .D(_0239_),
    .RESET_B(net23),
    .Q(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[23] ));
 sky130_fd_sc_hd__dfrtp_1 _4426_ (.CLK(clknet_leaf_0_user_clock2),
    .D(_0240_),
    .RESET_B(net12),
    .Q(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[24] ));
 sky130_fd_sc_hd__dfrtp_1 _4427_ (.CLK(clknet_leaf_2_user_clock2),
    .D(_0241_),
    .RESET_B(net24),
    .Q(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[25] ));
 sky130_fd_sc_hd__dfrtp_1 _4428_ (.CLK(clknet_leaf_0_user_clock2),
    .D(_0242_),
    .RESET_B(net13),
    .Q(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[26] ));
 sky130_fd_sc_hd__dfrtp_1 _4429_ (.CLK(clknet_leaf_0_user_clock2),
    .D(_0243_),
    .RESET_B(net14),
    .Q(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[27] ));
 sky130_fd_sc_hd__dfrtp_1 _4430_ (.CLK(clknet_leaf_0_user_clock2),
    .D(_0244_),
    .RESET_B(net11),
    .Q(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[28] ));
 sky130_fd_sc_hd__dfrtp_1 _4431_ (.CLK(clknet_leaf_1_user_clock2),
    .D(_0245_),
    .RESET_B(net17),
    .Q(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[29] ));
 sky130_fd_sc_hd__dfrtp_1 _4432_ (.CLK(clknet_leaf_2_user_clock2),
    .D(_0246_),
    .RESET_B(net18),
    .Q(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[30] ));
 sky130_fd_sc_hd__dfrtp_1 _4433_ (.CLK(clknet_leaf_2_user_clock2),
    .D(_0247_),
    .RESET_B(net24),
    .Q(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[31] ));
 sky130_fd_sc_hd__dfrtp_1 _4434_ (.CLK(clknet_leaf_0_user_clock2),
    .D(_0248_),
    .RESET_B(net11),
    .Q(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[32] ));
 sky130_fd_sc_hd__dfrtp_1 _4435_ (.CLK(clknet_leaf_2_user_clock2),
    .D(_0249_),
    .RESET_B(net16),
    .Q(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[33] ));
 sky130_fd_sc_hd__dfrtp_1 _4436_ (.CLK(clknet_leaf_37_user_clock2),
    .D(_0250_),
    .RESET_B(net11),
    .Q(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[34] ));
 sky130_fd_sc_hd__dfrtp_1 _4437_ (.CLK(clknet_leaf_37_user_clock2),
    .D(_0251_),
    .RESET_B(net11),
    .Q(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[35] ));
 sky130_fd_sc_hd__dfrtp_1 _4438_ (.CLK(clknet_leaf_37_user_clock2),
    .D(_0252_),
    .RESET_B(net12),
    .Q(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[36] ));
 sky130_fd_sc_hd__dfrtp_1 _4439_ (.CLK(clknet_leaf_37_user_clock2),
    .D(_0253_),
    .RESET_B(net18),
    .Q(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[37] ));
 sky130_fd_sc_hd__dfrtp_1 _4440_ (.CLK(clknet_leaf_34_user_clock2),
    .D(_0254_),
    .RESET_B(net23),
    .Q(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[38] ));
 sky130_fd_sc_hd__dfrtp_1 _4441_ (.CLK(clknet_leaf_34_user_clock2),
    .D(_0255_),
    .RESET_B(net25),
    .Q(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[39] ));
 sky130_fd_sc_hd__dfrtp_1 _4442_ (.CLK(clknet_leaf_0_user_clock2),
    .D(_0256_),
    .RESET_B(net11),
    .Q(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[40] ));
 sky130_fd_sc_hd__dfrtp_1 _4443_ (.CLK(clknet_leaf_2_user_clock2),
    .D(_0257_),
    .RESET_B(net23),
    .Q(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[41] ));
 sky130_fd_sc_hd__dfrtp_1 _4444_ (.CLK(clknet_leaf_37_user_clock2),
    .D(_0258_),
    .RESET_B(net11),
    .Q(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[42] ));
 sky130_fd_sc_hd__dfrtp_1 _4445_ (.CLK(clknet_leaf_37_user_clock2),
    .D(_0259_),
    .RESET_B(net12),
    .Q(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[43] ));
 sky130_fd_sc_hd__dfrtp_1 _4446_ (.CLK(clknet_leaf_37_user_clock2),
    .D(_0260_),
    .RESET_B(net12),
    .Q(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[44] ));
 sky130_fd_sc_hd__dfrtp_1 _4447_ (.CLK(clknet_leaf_34_user_clock2),
    .D(_0261_),
    .RESET_B(net18),
    .Q(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[45] ));
 sky130_fd_sc_hd__dfrtp_1 _4448_ (.CLK(clknet_leaf_36_user_clock2),
    .D(_0262_),
    .RESET_B(net23),
    .Q(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[46] ));
 sky130_fd_sc_hd__dfrtp_1 _4449_ (.CLK(clknet_leaf_34_user_clock2),
    .D(_0263_),
    .RESET_B(net25),
    .Q(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[47] ));
 sky130_fd_sc_hd__dfrtp_1 _4450_ (.CLK(clknet_leaf_0_user_clock2),
    .D(_0264_),
    .RESET_B(net12),
    .Q(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[48] ));
 sky130_fd_sc_hd__dfrtp_1 _4451_ (.CLK(clknet_leaf_2_user_clock2),
    .D(_0265_),
    .RESET_B(net23),
    .Q(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[49] ));
 sky130_fd_sc_hd__dfrtp_1 _4452_ (.CLK(clknet_leaf_0_user_clock2),
    .D(_0266_),
    .RESET_B(net11),
    .Q(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[50] ));
 sky130_fd_sc_hd__dfrtp_1 _4453_ (.CLK(clknet_leaf_0_user_clock2),
    .D(_0267_),
    .RESET_B(net12),
    .Q(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[51] ));
 sky130_fd_sc_hd__dfrtp_1 _4454_ (.CLK(clknet_leaf_0_user_clock2),
    .D(_0268_),
    .RESET_B(net11),
    .Q(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[52] ));
 sky130_fd_sc_hd__dfrtp_1 _4455_ (.CLK(clknet_leaf_37_user_clock2),
    .D(_0269_),
    .RESET_B(net16),
    .Q(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[53] ));
 sky130_fd_sc_hd__dfrtp_1 _4456_ (.CLK(clknet_leaf_2_user_clock2),
    .D(_0270_),
    .RESET_B(net18),
    .Q(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[54] ));
 sky130_fd_sc_hd__dfrtp_1 _4457_ (.CLK(clknet_leaf_33_user_clock2),
    .D(_0271_),
    .RESET_B(net23),
    .Q(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[55] ));
 sky130_fd_sc_hd__dfrtp_1 _4458_ (.CLK(clknet_leaf_0_user_clock2),
    .D(_0272_),
    .RESET_B(net12),
    .Q(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[56] ));
 sky130_fd_sc_hd__dfrtp_1 _4459_ (.CLK(clknet_leaf_33_user_clock2),
    .D(_0273_),
    .RESET_B(net23),
    .Q(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[57] ));
 sky130_fd_sc_hd__dfrtp_1 _4460_ (.CLK(clknet_leaf_37_user_clock2),
    .D(_0274_),
    .RESET_B(net11),
    .Q(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[58] ));
 sky130_fd_sc_hd__dfrtp_1 _4461_ (.CLK(clknet_leaf_0_user_clock2),
    .D(_0275_),
    .RESET_B(net12),
    .Q(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[59] ));
 sky130_fd_sc_hd__dfrtp_1 _4462_ (.CLK(clknet_leaf_0_user_clock2),
    .D(_0276_),
    .RESET_B(net15),
    .Q(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[60] ));
 sky130_fd_sc_hd__dfrtp_1 _4463_ (.CLK(clknet_leaf_37_user_clock2),
    .D(_0277_),
    .RESET_B(net16),
    .Q(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[61] ));
 sky130_fd_sc_hd__dfrtp_1 _4464_ (.CLK(clknet_leaf_33_user_clock2),
    .D(_0278_),
    .RESET_B(net23),
    .Q(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[62] ));
 sky130_fd_sc_hd__dfrtp_1 _4465_ (.CLK(clknet_leaf_33_user_clock2),
    .D(_0279_),
    .RESET_B(net23),
    .Q(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[63] ));
 sky130_fd_sc_hd__dfrtp_1 _4466_ (.CLK(clknet_leaf_37_user_clock2),
    .D(_0280_),
    .RESET_B(net16),
    .Q(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[64] ));
 sky130_fd_sc_hd__dfrtp_1 _4467_ (.CLK(clknet_leaf_2_user_clock2),
    .D(_0281_),
    .RESET_B(net16),
    .Q(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[65] ));
 sky130_fd_sc_hd__dfrtp_1 _4468_ (.CLK(clknet_leaf_37_user_clock2),
    .D(_0282_),
    .RESET_B(net16),
    .Q(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[66] ));
 sky130_fd_sc_hd__dfrtp_1 _4469_ (.CLK(clknet_leaf_37_user_clock2),
    .D(_0283_),
    .RESET_B(net12),
    .Q(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[67] ));
 sky130_fd_sc_hd__dfrtp_1 _4470_ (.CLK(clknet_leaf_37_user_clock2),
    .D(_0284_),
    .RESET_B(net16),
    .Q(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[68] ));
 sky130_fd_sc_hd__dfrtp_1 _4471_ (.CLK(clknet_leaf_37_user_clock2),
    .D(_0285_),
    .RESET_B(net16),
    .Q(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[69] ));
 sky130_fd_sc_hd__dfrtp_1 _4472_ (.CLK(clknet_leaf_2_user_clock2),
    .D(_0286_),
    .RESET_B(net16),
    .Q(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[70] ));
 sky130_fd_sc_hd__dfrtp_1 _4473_ (.CLK(clknet_leaf_2_user_clock2),
    .D(_0287_),
    .RESET_B(net25),
    .Q(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_fifo_q[71] ));
 sky130_fd_sc_hd__dfrtp_1 _4474_ (.CLK(clknet_leaf_34_user_clock2),
    .D(_0288_),
    .RESET_B(net26),
    .Q(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.delay_out_cnt_q[0] ));
 sky130_fd_sc_hd__dfrtp_1 _4475_ (.CLK(clknet_leaf_34_user_clock2),
    .D(_0289_),
    .RESET_B(net26),
    .Q(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.delay_out_cnt_q[1] ));
 sky130_fd_sc_hd__dfrtp_1 _4476_ (.CLK(clknet_leaf_20_user_clock2),
    .D(_0290_),
    .RESET_B(net46),
    .Q(\usb2uart.u_usb_cdc.bulk_in_valid ));
 sky130_fd_sc_hd__dfrtp_4 _4477_ (.CLK(clknet_leaf_34_user_clock2),
    .D(_0291_),
    .RESET_B(net26),
    .Q(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_first_q[0] ));
 sky130_fd_sc_hd__dfrtp_1 _4478_ (.CLK(clknet_leaf_34_user_clock2),
    .D(_0292_),
    .RESET_B(net26),
    .Q(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_first_q[1] ));
 sky130_fd_sc_hd__dfrtp_4 _4479_ (.CLK(clknet_leaf_33_user_clock2),
    .D(_0293_),
    .RESET_B(net26),
    .Q(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_first_q[2] ));
 sky130_fd_sc_hd__dfrtp_2 _4480_ (.CLK(clknet_leaf_33_user_clock2),
    .D(_0294_),
    .RESET_B(net26),
    .Q(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_first_q[3] ));
 sky130_fd_sc_hd__dfrtp_1 _4481_ (.CLK(clknet_leaf_33_user_clock2),
    .D(_0295_),
    .RESET_B(net26),
    .Q(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_full_o ));
 sky130_fd_sc_hd__dfrtp_1 _4482_ (.CLK(clknet_leaf_24_user_clock2),
    .D(_0296_),
    .RESET_B(net49),
    .Q(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_first_qq[0] ));
 sky130_fd_sc_hd__dfrtp_1 _4483_ (.CLK(clknet_leaf_24_user_clock2),
    .D(_0297_),
    .RESET_B(net49),
    .Q(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_first_qq[1] ));
 sky130_fd_sc_hd__dfrtp_1 _4484_ (.CLK(clknet_leaf_23_user_clock2),
    .D(_0298_),
    .RESET_B(net46),
    .Q(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_first_qq[2] ));
 sky130_fd_sc_hd__dfrtp_4 _4485_ (.CLK(clknet_leaf_22_user_clock2),
    .D(_0299_),
    .RESET_B(net37),
    .Q(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_first_qq[3] ));
 sky130_fd_sc_hd__dfrtp_1 _4486_ (.CLK(clknet_leaf_21_user_clock2),
    .D(_0038_),
    .RESET_B(net38),
    .Q(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_state_q ));
 sky130_fd_sc_hd__dfrtp_2 _4487_ (.CLK(clknet_leaf_21_user_clock2),
    .D(\usb2uart.u_usb_cdc.bulk_in_req ),
    .RESET_B(net46),
    .Q(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_req_q ));
 sky130_fd_sc_hd__dfrtp_1 _4488_ (.CLK(clknet_leaf_20_user_clock2),
    .D(_0300_),
    .RESET_B(net46),
    .Q(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_first_q[0] ));
 sky130_fd_sc_hd__dfrtp_1 _4489_ (.CLK(clknet_leaf_20_user_clock2),
    .D(_0301_),
    .RESET_B(net46),
    .Q(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_first_q[1] ));
 sky130_fd_sc_hd__dfrtp_1 _4490_ (.CLK(clknet_leaf_22_user_clock2),
    .D(_0302_),
    .RESET_B(net37),
    .Q(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_first_q[2] ));
 sky130_fd_sc_hd__dfrtp_2 _4491_ (.CLK(clknet_leaf_21_user_clock2),
    .D(_0303_),
    .RESET_B(net37),
    .Q(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_first_q[3] ));
 sky130_fd_sc_hd__dfrtp_1 _4492_ (.CLK(clknet_leaf_32_user_clock2),
    .D(_0304_),
    .RESET_B(net33),
    .Q(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.delay_in_cnt_q[0] ));
 sky130_fd_sc_hd__dfrtp_1 _4493_ (.CLK(clknet_leaf_32_user_clock2),
    .D(_0305_),
    .RESET_B(net33),
    .Q(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.delay_in_cnt_q[1] ));
 sky130_fd_sc_hd__dfxtp_1 _4494_ (.CLK(clknet_leaf_36_user_clock2),
    .D(_0306_),
    .Q(\usb2uart.u_uart.uart_tx_inst.data_reg[0] ));
 sky130_fd_sc_hd__dfxtp_1 _4495_ (.CLK(clknet_leaf_36_user_clock2),
    .D(_0307_),
    .Q(\usb2uart.u_uart.uart_tx_inst.data_reg[1] ));
 sky130_fd_sc_hd__dfxtp_1 _4496_ (.CLK(clknet_leaf_36_user_clock2),
    .D(_0308_),
    .Q(\usb2uart.u_uart.uart_tx_inst.data_reg[2] ));
 sky130_fd_sc_hd__dfxtp_1 _4497_ (.CLK(clknet_leaf_37_user_clock2),
    .D(_0309_),
    .Q(\usb2uart.u_uart.uart_tx_inst.data_reg[3] ));
 sky130_fd_sc_hd__dfxtp_1 _4498_ (.CLK(clknet_leaf_37_user_clock2),
    .D(_0310_),
    .Q(\usb2uart.u_uart.uart_tx_inst.data_reg[4] ));
 sky130_fd_sc_hd__dfxtp_1 _4499_ (.CLK(clknet_leaf_36_user_clock2),
    .D(_0311_),
    .Q(\usb2uart.u_uart.uart_tx_inst.data_reg[5] ));
 sky130_fd_sc_hd__dfxtp_1 _4500_ (.CLK(clknet_leaf_36_user_clock2),
    .D(_0312_),
    .Q(\usb2uart.u_uart.uart_tx_inst.data_reg[6] ));
 sky130_fd_sc_hd__dfxtp_1 _4501_ (.CLK(clknet_leaf_36_user_clock2),
    .D(_0313_),
    .Q(\usb2uart.u_uart.uart_tx_inst.data_reg[7] ));
 sky130_fd_sc_hd__dfxtp_1 _4502_ (.CLK(clknet_leaf_34_user_clock2),
    .D(_0314_),
    .Q(\usb2uart.u_uart.uart_tx_inst.data_reg[8] ));
 sky130_fd_sc_hd__dfrtp_1 _4503_ (.CLK(clknet_leaf_26_user_clock2),
    .D(_0315_),
    .RESET_B(net48),
    .Q(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[0] ));
 sky130_fd_sc_hd__dfrtp_1 _4504_ (.CLK(clknet_leaf_26_user_clock2),
    .D(_0316_),
    .RESET_B(net47),
    .Q(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[1] ));
 sky130_fd_sc_hd__dfrtp_1 _4505_ (.CLK(clknet_leaf_26_user_clock2),
    .D(_0317_),
    .RESET_B(net45),
    .Q(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[2] ));
 sky130_fd_sc_hd__dfrtp_1 _4506_ (.CLK(clknet_leaf_27_user_clock2),
    .D(_0318_),
    .RESET_B(net44),
    .Q(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[3] ));
 sky130_fd_sc_hd__dfrtp_1 _4507_ (.CLK(clknet_leaf_27_user_clock2),
    .D(_0319_),
    .RESET_B(net44),
    .Q(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[4] ));
 sky130_fd_sc_hd__dfrtp_1 _4508_ (.CLK(clknet_leaf_26_user_clock2),
    .D(_0320_),
    .RESET_B(net45),
    .Q(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[5] ));
 sky130_fd_sc_hd__dfrtp_1 _4509_ (.CLK(clknet_leaf_24_user_clock2),
    .D(_0321_),
    .RESET_B(net47),
    .Q(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[6] ));
 sky130_fd_sc_hd__dfrtp_1 _4510_ (.CLK(clknet_leaf_27_user_clock2),
    .D(_0322_),
    .RESET_B(net44),
    .Q(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[7] ));
 sky130_fd_sc_hd__dfrtp_1 _4511_ (.CLK(clknet_leaf_25_user_clock2),
    .D(_0323_),
    .RESET_B(net48),
    .Q(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[8] ));
 sky130_fd_sc_hd__dfrtp_1 _4512_ (.CLK(clknet_leaf_26_user_clock2),
    .D(_0324_),
    .RESET_B(net47),
    .Q(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[9] ));
 sky130_fd_sc_hd__dfrtp_1 _4513_ (.CLK(clknet_leaf_26_user_clock2),
    .D(_0325_),
    .RESET_B(net47),
    .Q(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[10] ));
 sky130_fd_sc_hd__dfrtp_1 _4514_ (.CLK(clknet_leaf_26_user_clock2),
    .D(_0326_),
    .RESET_B(net45),
    .Q(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[11] ));
 sky130_fd_sc_hd__dfrtp_1 _4515_ (.CLK(clknet_leaf_26_user_clock2),
    .D(_0327_),
    .RESET_B(net44),
    .Q(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[12] ));
 sky130_fd_sc_hd__dfrtp_1 _4516_ (.CLK(clknet_leaf_26_user_clock2),
    .D(_0328_),
    .RESET_B(net45),
    .Q(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[13] ));
 sky130_fd_sc_hd__dfrtp_1 _4517_ (.CLK(clknet_leaf_25_user_clock2),
    .D(_0329_),
    .RESET_B(net48),
    .Q(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[14] ));
 sky130_fd_sc_hd__dfrtp_1 _4518_ (.CLK(clknet_leaf_26_user_clock2),
    .D(_0330_),
    .RESET_B(net45),
    .Q(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[15] ));
 sky130_fd_sc_hd__dfrtp_1 _4519_ (.CLK(clknet_leaf_25_user_clock2),
    .D(_0331_),
    .RESET_B(net48),
    .Q(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[16] ));
 sky130_fd_sc_hd__dfrtp_1 _4520_ (.CLK(clknet_leaf_25_user_clock2),
    .D(_0332_),
    .RESET_B(net45),
    .Q(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[17] ));
 sky130_fd_sc_hd__dfrtp_1 _4521_ (.CLK(clknet_leaf_22_user_clock2),
    .D(_0333_),
    .RESET_B(net34),
    .Q(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[18] ));
 sky130_fd_sc_hd__dfrtp_1 _4522_ (.CLK(clknet_leaf_31_user_clock2),
    .D(_0334_),
    .RESET_B(net35),
    .Q(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[19] ));
 sky130_fd_sc_hd__dfrtp_1 _4523_ (.CLK(clknet_leaf_31_user_clock2),
    .D(_0335_),
    .RESET_B(net33),
    .Q(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[20] ));
 sky130_fd_sc_hd__dfrtp_1 _4524_ (.CLK(clknet_leaf_31_user_clock2),
    .D(_0336_),
    .RESET_B(net33),
    .Q(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[21] ));
 sky130_fd_sc_hd__dfrtp_1 _4525_ (.CLK(clknet_leaf_24_user_clock2),
    .D(_0337_),
    .RESET_B(net49),
    .Q(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[22] ));
 sky130_fd_sc_hd__dfrtp_1 _4526_ (.CLK(clknet_leaf_31_user_clock2),
    .D(_0338_),
    .RESET_B(net34),
    .Q(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[23] ));
 sky130_fd_sc_hd__dfrtp_1 _4527_ (.CLK(clknet_leaf_25_user_clock2),
    .D(_0339_),
    .RESET_B(net47),
    .Q(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[24] ));
 sky130_fd_sc_hd__dfrtp_1 _4528_ (.CLK(clknet_leaf_25_user_clock2),
    .D(_0340_),
    .RESET_B(net47),
    .Q(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[25] ));
 sky130_fd_sc_hd__dfrtp_1 _4529_ (.CLK(clknet_leaf_22_user_clock2),
    .D(_0341_),
    .RESET_B(net37),
    .Q(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[26] ));
 sky130_fd_sc_hd__dfrtp_1 _4530_ (.CLK(clknet_leaf_30_user_clock2),
    .D(_0342_),
    .RESET_B(net35),
    .Q(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[27] ));
 sky130_fd_sc_hd__dfrtp_1 _4531_ (.CLK(clknet_leaf_32_user_clock2),
    .D(_0343_),
    .RESET_B(net33),
    .Q(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[28] ));
 sky130_fd_sc_hd__dfrtp_1 _4532_ (.CLK(clknet_leaf_31_user_clock2),
    .D(_0344_),
    .RESET_B(net33),
    .Q(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[29] ));
 sky130_fd_sc_hd__dfrtp_1 _4533_ (.CLK(clknet_leaf_24_user_clock2),
    .D(_0345_),
    .RESET_B(net53),
    .Q(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[30] ));
 sky130_fd_sc_hd__dfrtp_1 _4534_ (.CLK(clknet_leaf_31_user_clock2),
    .D(_0346_),
    .RESET_B(net33),
    .Q(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[31] ));
 sky130_fd_sc_hd__dfrtp_1 _4535_ (.CLK(clknet_leaf_25_user_clock2),
    .D(_0347_),
    .RESET_B(net48),
    .Q(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[32] ));
 sky130_fd_sc_hd__dfrtp_1 _4536_ (.CLK(clknet_leaf_26_user_clock2),
    .D(_0348_),
    .RESET_B(net45),
    .Q(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[33] ));
 sky130_fd_sc_hd__dfrtp_1 _4537_ (.CLK(clknet_leaf_22_user_clock2),
    .D(_0349_),
    .RESET_B(net38),
    .Q(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[34] ));
 sky130_fd_sc_hd__dfrtp_1 _4538_ (.CLK(clknet_leaf_30_user_clock2),
    .D(_0350_),
    .RESET_B(net35),
    .Q(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[35] ));
 sky130_fd_sc_hd__dfrtp_1 _4539_ (.CLK(clknet_leaf_31_user_clock2),
    .D(_0351_),
    .RESET_B(net35),
    .Q(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[36] ));
 sky130_fd_sc_hd__dfrtp_1 _4540_ (.CLK(clknet_leaf_31_user_clock2),
    .D(_0352_),
    .RESET_B(net36),
    .Q(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[37] ));
 sky130_fd_sc_hd__dfrtp_1 _4541_ (.CLK(clknet_leaf_24_user_clock2),
    .D(_0353_),
    .RESET_B(net49),
    .Q(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[38] ));
 sky130_fd_sc_hd__dfrtp_1 _4542_ (.CLK(clknet_leaf_31_user_clock2),
    .D(_0354_),
    .RESET_B(net35),
    .Q(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[39] ));
 sky130_fd_sc_hd__dfrtp_1 _4543_ (.CLK(clknet_leaf_25_user_clock2),
    .D(_0355_),
    .RESET_B(net48),
    .Q(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[40] ));
 sky130_fd_sc_hd__dfrtp_1 _4544_ (.CLK(clknet_leaf_25_user_clock2),
    .D(_0356_),
    .RESET_B(net47),
    .Q(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[41] ));
 sky130_fd_sc_hd__dfrtp_1 _4545_ (.CLK(clknet_leaf_31_user_clock2),
    .D(_0357_),
    .RESET_B(net36),
    .Q(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[42] ));
 sky130_fd_sc_hd__dfrtp_1 _4546_ (.CLK(clknet_leaf_27_user_clock2),
    .D(_0358_),
    .RESET_B(net36),
    .Q(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[43] ));
 sky130_fd_sc_hd__dfrtp_1 _4547_ (.CLK(clknet_leaf_31_user_clock2),
    .D(_0359_),
    .RESET_B(net36),
    .Q(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[44] ));
 sky130_fd_sc_hd__dfrtp_1 _4548_ (.CLK(clknet_leaf_31_user_clock2),
    .D(_0360_),
    .RESET_B(net36),
    .Q(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[45] ));
 sky130_fd_sc_hd__dfrtp_1 _4549_ (.CLK(clknet_leaf_25_user_clock2),
    .D(_0361_),
    .RESET_B(net48),
    .Q(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[46] ));
 sky130_fd_sc_hd__dfrtp_1 _4550_ (.CLK(clknet_leaf_27_user_clock2),
    .D(_0362_),
    .RESET_B(net36),
    .Q(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[47] ));
 sky130_fd_sc_hd__dfrtp_1 _4551_ (.CLK(clknet_leaf_24_user_clock2),
    .D(_0363_),
    .RESET_B(net47),
    .Q(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[48] ));
 sky130_fd_sc_hd__dfrtp_1 _4552_ (.CLK(clknet_leaf_23_user_clock2),
    .D(_0364_),
    .RESET_B(net45),
    .Q(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[49] ));
 sky130_fd_sc_hd__dfrtp_1 _4553_ (.CLK(clknet_leaf_23_user_clock2),
    .D(_0365_),
    .RESET_B(net37),
    .Q(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[50] ));
 sky130_fd_sc_hd__dfrtp_1 _4554_ (.CLK(clknet_leaf_31_user_clock2),
    .D(_0366_),
    .RESET_B(net35),
    .Q(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[51] ));
 sky130_fd_sc_hd__dfrtp_1 _4555_ (.CLK(clknet_leaf_31_user_clock2),
    .D(_0367_),
    .RESET_B(net35),
    .Q(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[52] ));
 sky130_fd_sc_hd__dfrtp_1 _4556_ (.CLK(clknet_leaf_22_user_clock2),
    .D(_0368_),
    .RESET_B(net36),
    .Q(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[53] ));
 sky130_fd_sc_hd__dfrtp_1 _4557_ (.CLK(clknet_leaf_24_user_clock2),
    .D(_0369_),
    .RESET_B(net49),
    .Q(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[54] ));
 sky130_fd_sc_hd__dfrtp_1 _4558_ (.CLK(clknet_leaf_31_user_clock2),
    .D(_0370_),
    .RESET_B(net35),
    .Q(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[55] ));
 sky130_fd_sc_hd__dfrtp_1 _4559_ (.CLK(clknet_leaf_25_user_clock2),
    .D(_0371_),
    .RESET_B(net47),
    .Q(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[56] ));
 sky130_fd_sc_hd__dfrtp_1 _4560_ (.CLK(clknet_leaf_23_user_clock2),
    .D(_0372_),
    .RESET_B(net44),
    .Q(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[57] ));
 sky130_fd_sc_hd__dfrtp_1 _4561_ (.CLK(clknet_leaf_23_user_clock2),
    .D(_0373_),
    .RESET_B(net46),
    .Q(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[58] ));
 sky130_fd_sc_hd__dfrtp_1 _4562_ (.CLK(clknet_leaf_23_user_clock2),
    .D(_0374_),
    .RESET_B(net44),
    .Q(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[59] ));
 sky130_fd_sc_hd__dfrtp_1 _4563_ (.CLK(clknet_leaf_23_user_clock2),
    .D(_0375_),
    .RESET_B(net44),
    .Q(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[60] ));
 sky130_fd_sc_hd__dfrtp_1 _4564_ (.CLK(clknet_leaf_23_user_clock2),
    .D(_0376_),
    .RESET_B(net44),
    .Q(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[61] ));
 sky130_fd_sc_hd__dfrtp_1 _4565_ (.CLK(clknet_leaf_24_user_clock2),
    .D(_0377_),
    .RESET_B(net53),
    .Q(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[62] ));
 sky130_fd_sc_hd__dfrtp_1 _4566_ (.CLK(clknet_leaf_23_user_clock2),
    .D(_0378_),
    .RESET_B(net44),
    .Q(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[63] ));
 sky130_fd_sc_hd__dfrtp_1 _4567_ (.CLK(clknet_leaf_25_user_clock2),
    .D(_0379_),
    .RESET_B(net47),
    .Q(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[64] ));
 sky130_fd_sc_hd__dfrtp_1 _4568_ (.CLK(clknet_leaf_23_user_clock2),
    .D(_0380_),
    .RESET_B(net44),
    .Q(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[65] ));
 sky130_fd_sc_hd__dfrtp_1 _4569_ (.CLK(clknet_leaf_22_user_clock2),
    .D(_0381_),
    .RESET_B(net37),
    .Q(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[66] ));
 sky130_fd_sc_hd__dfrtp_1 _4570_ (.CLK(clknet_leaf_22_user_clock2),
    .D(_0382_),
    .RESET_B(net37),
    .Q(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[67] ));
 sky130_fd_sc_hd__dfrtp_1 _4571_ (.CLK(clknet_leaf_22_user_clock2),
    .D(_0383_),
    .RESET_B(net35),
    .Q(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[68] ));
 sky130_fd_sc_hd__dfrtp_1 _4572_ (.CLK(clknet_leaf_31_user_clock2),
    .D(_0384_),
    .RESET_B(net35),
    .Q(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[69] ));
 sky130_fd_sc_hd__dfrtp_1 _4573_ (.CLK(clknet_leaf_23_user_clock2),
    .D(_0385_),
    .RESET_B(net46),
    .Q(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[70] ));
 sky130_fd_sc_hd__dfrtp_1 _4574_ (.CLK(clknet_leaf_22_user_clock2),
    .D(_0386_),
    .RESET_B(net37),
    .Q(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_fifo_q[71] ));
 sky130_fd_sc_hd__dfrtp_4 _4575_ (.CLK(clknet_leaf_24_user_clock2),
    .D(_0387_),
    .RESET_B(net49),
    .Q(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_last_q[0] ));
 sky130_fd_sc_hd__dfrtp_4 _4576_ (.CLK(clknet_leaf_24_user_clock2),
    .D(_0388_),
    .RESET_B(net49),
    .Q(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_last_q[1] ));
 sky130_fd_sc_hd__dfrtp_4 _4577_ (.CLK(clknet_leaf_24_user_clock2),
    .D(_0389_),
    .RESET_B(net49),
    .Q(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_last_q[2] ));
 sky130_fd_sc_hd__dfrtp_4 _4578_ (.CLK(clknet_leaf_24_user_clock2),
    .D(_0390_),
    .RESET_B(net46),
    .Q(\usb2uart.u_usb_cdc.u_bulk_endp.u_in_fifo.in_last_q[3] ));
 sky130_fd_sc_hd__dfxtp_1 _4579_ (.CLK(clknet_leaf_34_user_clock2),
    .D(_0391_),
    .Q(\usb2uart.u_uart.uart_tx_inst.prescale_reg[0] ));
 sky130_fd_sc_hd__dfxtp_1 _4580_ (.CLK(clknet_leaf_35_user_clock2),
    .D(_0392_),
    .Q(\usb2uart.u_uart.uart_tx_inst.prescale_reg[1] ));
 sky130_fd_sc_hd__dfxtp_1 _4581_ (.CLK(clknet_leaf_35_user_clock2),
    .D(_0393_),
    .Q(\usb2uart.u_uart.uart_tx_inst.prescale_reg[2] ));
 sky130_fd_sc_hd__dfxtp_1 _4582_ (.CLK(clknet_leaf_35_user_clock2),
    .D(_0394_),
    .Q(\usb2uart.u_uart.uart_tx_inst.prescale_reg[3] ));
 sky130_fd_sc_hd__dfxtp_1 _4583_ (.CLK(clknet_leaf_35_user_clock2),
    .D(_0395_),
    .Q(\usb2uart.u_uart.uart_tx_inst.prescale_reg[4] ));
 sky130_fd_sc_hd__dfxtp_1 _4584_ (.CLK(clknet_leaf_35_user_clock2),
    .D(_0396_),
    .Q(\usb2uart.u_uart.uart_tx_inst.prescale_reg[5] ));
 sky130_fd_sc_hd__dfxtp_1 _4585_ (.CLK(clknet_leaf_35_user_clock2),
    .D(_0397_),
    .Q(\usb2uart.u_uart.uart_tx_inst.prescale_reg[6] ));
 sky130_fd_sc_hd__dfxtp_1 _4586_ (.CLK(clknet_leaf_35_user_clock2),
    .D(_0398_),
    .Q(\usb2uart.u_uart.uart_tx_inst.prescale_reg[7] ));
 sky130_fd_sc_hd__dfxtp_1 _4587_ (.CLK(clknet_leaf_35_user_clock2),
    .D(_0399_),
    .Q(\usb2uart.u_uart.uart_tx_inst.prescale_reg[8] ));
 sky130_fd_sc_hd__dfxtp_1 _4588_ (.CLK(clknet_leaf_35_user_clock2),
    .D(_0400_),
    .Q(\usb2uart.u_uart.uart_tx_inst.prescale_reg[9] ));
 sky130_fd_sc_hd__dfxtp_1 _4589_ (.CLK(clknet_leaf_35_user_clock2),
    .D(_0401_),
    .Q(\usb2uart.u_uart.uart_tx_inst.prescale_reg[10] ));
 sky130_fd_sc_hd__dfxtp_1 _4590_ (.CLK(clknet_leaf_35_user_clock2),
    .D(_0402_),
    .Q(\usb2uart.u_uart.uart_tx_inst.prescale_reg[11] ));
 sky130_fd_sc_hd__dfxtp_1 _4591_ (.CLK(clknet_leaf_35_user_clock2),
    .D(_0403_),
    .Q(\usb2uart.u_uart.uart_tx_inst.prescale_reg[12] ));
 sky130_fd_sc_hd__dfxtp_1 _4592_ (.CLK(clknet_leaf_35_user_clock2),
    .D(_0404_),
    .Q(\usb2uart.u_uart.uart_tx_inst.prescale_reg[13] ));
 sky130_fd_sc_hd__dfxtp_1 _4593_ (.CLK(clknet_leaf_35_user_clock2),
    .D(_0405_),
    .Q(\usb2uart.u_uart.uart_tx_inst.prescale_reg[14] ));
 sky130_fd_sc_hd__dfxtp_1 _4594_ (.CLK(clknet_leaf_30_user_clock2),
    .D(_0406_),
    .Q(\usb2uart.u_uart.uart_tx_inst.prescale_reg[15] ));
 sky130_fd_sc_hd__dfxtp_1 _4595_ (.CLK(clknet_leaf_29_user_clock2),
    .D(_0407_),
    .Q(\usb2uart.u_uart.uart_tx_inst.prescale_reg[16] ));
 sky130_fd_sc_hd__dfxtp_1 _4596_ (.CLK(clknet_leaf_35_user_clock2),
    .D(_0408_),
    .Q(\usb2uart.u_uart.uart_tx_inst.prescale_reg[17] ));
 sky130_fd_sc_hd__dfxtp_1 _4597_ (.CLK(clknet_leaf_35_user_clock2),
    .D(_0409_),
    .Q(\usb2uart.u_uart.uart_tx_inst.prescale_reg[18] ));
 sky130_fd_sc_hd__dfxtp_1 _4598_ (.CLK(clknet_leaf_34_user_clock2),
    .D(_0410_),
    .Q(\usb2uart.u_uart.uart_tx_inst.bit_cnt[0] ));
 sky130_fd_sc_hd__dfxtp_1 _4599_ (.CLK(clknet_leaf_34_user_clock2),
    .D(_0411_),
    .Q(\usb2uart.u_uart.uart_tx_inst.bit_cnt[1] ));
 sky130_fd_sc_hd__dfxtp_1 _4600_ (.CLK(clknet_leaf_34_user_clock2),
    .D(_0412_),
    .Q(\usb2uart.u_uart.uart_tx_inst.bit_cnt[2] ));
 sky130_fd_sc_hd__dfxtp_1 _4601_ (.CLK(clknet_leaf_30_user_clock2),
    .D(_0413_),
    .Q(\usb2uart.u_uart.uart_tx_inst.bit_cnt[3] ));
 sky130_fd_sc_hd__dfxtp_1 _4602_ (.CLK(clknet_leaf_34_user_clock2),
    .D(_0414_),
    .Q(\usb2uart.u_uart.uart_tx_inst.s_axis_tready_reg ));
 sky130_fd_sc_hd__dfxtp_2 _4603_ (.CLK(clknet_leaf_34_user_clock2),
    .D(_0415_),
    .Q(net10));
 sky130_fd_sc_hd__dfxtp_1 _4604_ (.CLK(clknet_leaf_30_user_clock2),
    .D(_0416_),
    .Q(\usb2uart.u_uart.uart_rx_inst.m_axis_tvalid_reg ));
 sky130_fd_sc_hd__dfrtp_1 _4605_ (.CLK(clknet_leaf_12_user_clock2),
    .D(_0417_),
    .RESET_B(net29),
    .Q(\usb2uart.u_usb_cdc.u_sie.datain_toggle_q[1] ));
 sky130_fd_sc_hd__dfxtp_2 _4606_ (.CLK(clknet_leaf_27_user_clock2),
    .D(_0418_),
    .Q(\usb2uart.u_uart.uart_rx_inst.m_axis_tdata_reg[0] ));
 sky130_fd_sc_hd__dfxtp_2 _4607_ (.CLK(clknet_leaf_27_user_clock2),
    .D(_0419_),
    .Q(\usb2uart.u_uart.uart_rx_inst.m_axis_tdata_reg[1] ));
 sky130_fd_sc_hd__dfxtp_2 _4608_ (.CLK(clknet_leaf_30_user_clock2),
    .D(_0420_),
    .Q(\usb2uart.u_uart.uart_rx_inst.m_axis_tdata_reg[2] ));
 sky130_fd_sc_hd__dfxtp_1 _4609_ (.CLK(clknet_leaf_30_user_clock2),
    .D(_0421_),
    .Q(\usb2uart.u_uart.uart_rx_inst.m_axis_tdata_reg[3] ));
 sky130_fd_sc_hd__dfxtp_2 _4610_ (.CLK(clknet_leaf_30_user_clock2),
    .D(_0422_),
    .Q(\usb2uart.u_uart.uart_rx_inst.m_axis_tdata_reg[4] ));
 sky130_fd_sc_hd__dfxtp_2 _4611_ (.CLK(clknet_leaf_30_user_clock2),
    .D(_0423_),
    .Q(\usb2uart.u_uart.uart_rx_inst.m_axis_tdata_reg[5] ));
 sky130_fd_sc_hd__dfxtp_2 _4612_ (.CLK(clknet_leaf_30_user_clock2),
    .D(_0424_),
    .Q(\usb2uart.u_uart.uart_rx_inst.m_axis_tdata_reg[6] ));
 sky130_fd_sc_hd__dfxtp_2 _4613_ (.CLK(clknet_leaf_30_user_clock2),
    .D(_0425_),
    .Q(\usb2uart.u_uart.uart_rx_inst.m_axis_tdata_reg[7] ));
 sky130_fd_sc_hd__dfxtp_2 _4614_ (.CLK(clknet_leaf_30_user_clock2),
    .D(_0426_),
    .Q(\usb2uart.u_uart.uart_rx_inst.rxd_reg ));
 sky130_fd_sc_hd__dfxtp_1 _4615_ (.CLK(clknet_leaf_27_user_clock2),
    .D(_0427_),
    .Q(\usb2uart.u_uart.uart_rx_inst.prescale_reg[0] ));
 sky130_fd_sc_hd__dfxtp_1 _4616_ (.CLK(clknet_leaf_28_user_clock2),
    .D(_0428_),
    .Q(\usb2uart.u_uart.uart_rx_inst.prescale_reg[1] ));
 sky130_fd_sc_hd__dfxtp_1 _4617_ (.CLK(clknet_leaf_27_user_clock2),
    .D(_0429_),
    .Q(\usb2uart.u_uart.uart_rx_inst.prescale_reg[2] ));
 sky130_fd_sc_hd__dfxtp_1 _4618_ (.CLK(clknet_leaf_28_user_clock2),
    .D(_0430_),
    .Q(\usb2uart.u_uart.uart_rx_inst.prescale_reg[3] ));
 sky130_fd_sc_hd__dfxtp_1 _4619_ (.CLK(clknet_leaf_28_user_clock2),
    .D(_0431_),
    .Q(\usb2uart.u_uart.uart_rx_inst.prescale_reg[4] ));
 sky130_fd_sc_hd__dfxtp_1 _4620_ (.CLK(clknet_leaf_27_user_clock2),
    .D(_0432_),
    .Q(\usb2uart.u_uart.uart_rx_inst.prescale_reg[5] ));
 sky130_fd_sc_hd__dfxtp_1 _4621_ (.CLK(clknet_leaf_28_user_clock2),
    .D(_0433_),
    .Q(\usb2uart.u_uart.uart_rx_inst.prescale_reg[6] ));
 sky130_fd_sc_hd__dfxtp_1 _4622_ (.CLK(clknet_leaf_28_user_clock2),
    .D(_0434_),
    .Q(\usb2uart.u_uart.uart_rx_inst.prescale_reg[7] ));
 sky130_fd_sc_hd__dfxtp_1 _4623_ (.CLK(clknet_leaf_28_user_clock2),
    .D(_0435_),
    .Q(\usb2uart.u_uart.uart_rx_inst.prescale_reg[8] ));
 sky130_fd_sc_hd__dfxtp_1 _4624_ (.CLK(clknet_leaf_28_user_clock2),
    .D(_0436_),
    .Q(\usb2uart.u_uart.uart_rx_inst.prescale_reg[9] ));
 sky130_fd_sc_hd__dfxtp_1 _4625_ (.CLK(clknet_leaf_28_user_clock2),
    .D(_0437_),
    .Q(\usb2uart.u_uart.uart_rx_inst.prescale_reg[10] ));
 sky130_fd_sc_hd__dfxtp_1 _4626_ (.CLK(clknet_leaf_29_user_clock2),
    .D(_0438_),
    .Q(\usb2uart.u_uart.uart_rx_inst.prescale_reg[11] ));
 sky130_fd_sc_hd__dfxtp_1 _4627_ (.CLK(clknet_leaf_28_user_clock2),
    .D(_0439_),
    .Q(\usb2uart.u_uart.uart_rx_inst.prescale_reg[12] ));
 sky130_fd_sc_hd__dfxtp_1 _4628_ (.CLK(clknet_leaf_29_user_clock2),
    .D(_0440_),
    .Q(\usb2uart.u_uart.uart_rx_inst.prescale_reg[13] ));
 sky130_fd_sc_hd__dfxtp_1 _4629_ (.CLK(clknet_leaf_29_user_clock2),
    .D(_0441_),
    .Q(\usb2uart.u_uart.uart_rx_inst.prescale_reg[14] ));
 sky130_fd_sc_hd__dfxtp_1 _4630_ (.CLK(clknet_leaf_29_user_clock2),
    .D(_0442_),
    .Q(\usb2uart.u_uart.uart_rx_inst.prescale_reg[15] ));
 sky130_fd_sc_hd__dfxtp_1 _4631_ (.CLK(clknet_leaf_29_user_clock2),
    .D(_0443_),
    .Q(\usb2uart.u_uart.uart_rx_inst.prescale_reg[16] ));
 sky130_fd_sc_hd__dfxtp_1 _4632_ (.CLK(clknet_leaf_28_user_clock2),
    .D(_0444_),
    .Q(\usb2uart.u_uart.uart_rx_inst.prescale_reg[17] ));
 sky130_fd_sc_hd__dfxtp_1 _4633_ (.CLK(clknet_leaf_29_user_clock2),
    .D(_0445_),
    .Q(\usb2uart.u_uart.uart_rx_inst.prescale_reg[18] ));
 sky130_fd_sc_hd__dfxtp_1 _4634_ (.CLK(clknet_leaf_30_user_clock2),
    .D(_0446_),
    .Q(\usb2uart.u_uart.uart_rx_inst.bit_cnt[0] ));
 sky130_fd_sc_hd__dfxtp_1 _4635_ (.CLK(clknet_leaf_29_user_clock2),
    .D(_0447_),
    .Q(\usb2uart.u_uart.uart_rx_inst.bit_cnt[1] ));
 sky130_fd_sc_hd__dfxtp_1 _4636_ (.CLK(clknet_leaf_29_user_clock2),
    .D(_0448_),
    .Q(\usb2uart.u_uart.uart_rx_inst.bit_cnt[2] ));
 sky130_fd_sc_hd__dfxtp_1 _4637_ (.CLK(clknet_leaf_29_user_clock2),
    .D(_0449_),
    .Q(\usb2uart.u_uart.uart_rx_inst.bit_cnt[3] ));
 sky130_fd_sc_hd__conb_1 user_proj_example_264 (.HI(net264));
 sky130_fd_sc_hd__conb_1 user_proj_example_265 (.HI(net265));
 sky130_fd_sc_hd__conb_1 user_proj_example_266 (.HI(net266));
 sky130_fd_sc_hd__conb_1 user_proj_example_267 (.HI(net267));
 sky130_fd_sc_hd__conb_1 user_proj_example_268 (.HI(net268));
 sky130_fd_sc_hd__conb_1 user_proj_example_269 (.HI(net269));
 sky130_fd_sc_hd__conb_1 user_proj_example_270 (.HI(net270));
 sky130_fd_sc_hd__conb_1 user_proj_example_271 (.HI(net271));
 sky130_fd_sc_hd__conb_1 user_proj_example_272 (.HI(net272));
 sky130_fd_sc_hd__conb_1 user_proj_example_273 (.HI(net273));
 sky130_fd_sc_hd__conb_1 user_proj_example_274 (.HI(net274));
 sky130_fd_sc_hd__conb_1 user_proj_example_275 (.HI(net275));
 sky130_fd_sc_hd__conb_1 user_proj_example_276 (.HI(net276));
 sky130_fd_sc_hd__conb_1 user_proj_example_277 (.HI(net277));
 sky130_fd_sc_hd__conb_1 user_proj_example_278 (.HI(net278));
 sky130_fd_sc_hd__conb_1 user_proj_example_279 (.HI(net279));
 sky130_fd_sc_hd__conb_1 user_proj_example_280 (.HI(net280));
 sky130_fd_sc_hd__conb_1 user_proj_example_281 (.HI(net281));
 sky130_fd_sc_hd__conb_1 user_proj_example_282 (.HI(net282));
 sky130_fd_sc_hd__conb_1 user_proj_example_283 (.HI(net283));
 sky130_fd_sc_hd__conb_1 user_proj_example_284 (.HI(net284));
 sky130_fd_sc_hd__conb_1 user_proj_example_285 (.HI(net285));
 sky130_fd_sc_hd__conb_1 user_proj_example_286 (.HI(net286));
 sky130_fd_sc_hd__conb_1 user_proj_example_287 (.HI(net287));
 sky130_fd_sc_hd__conb_1 user_proj_example_288 (.HI(net288));
 sky130_fd_sc_hd__conb_1 user_proj_example_289 (.HI(net289));
 sky130_fd_sc_hd__conb_1 user_proj_example_290 (.HI(net290));
 sky130_fd_sc_hd__conb_1 user_proj_example_291 (.HI(net291));
 sky130_fd_sc_hd__conb_1 user_proj_example_292 (.HI(net292));
 sky130_fd_sc_hd__conb_1 user_proj_example_293 (.HI(net293));
 sky130_fd_sc_hd__conb_1 user_proj_example_294 (.HI(net294));
 sky130_fd_sc_hd__conb_1 user_proj_example_295 (.HI(net295));
 sky130_fd_sc_hd__conb_1 user_proj_example_296 (.HI(net296));
 sky130_fd_sc_hd__conb_1 user_proj_example_297 (.HI(net297));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_0_user_clock2 (.A(clknet_2_0__leaf_user_clock2),
    .X(clknet_leaf_0_user_clock2));
 sky130_fd_sc_hd__conb_1 user_proj_example_64 (.LO(net64));
 sky130_fd_sc_hd__conb_1 user_proj_example_65 (.LO(net65));
 sky130_fd_sc_hd__conb_1 user_proj_example_66 (.LO(net66));
 sky130_fd_sc_hd__conb_1 user_proj_example_67 (.LO(net67));
 sky130_fd_sc_hd__conb_1 user_proj_example_68 (.LO(net68));
 sky130_fd_sc_hd__conb_1 user_proj_example_69 (.LO(net69));
 sky130_fd_sc_hd__conb_1 user_proj_example_70 (.LO(net70));
 sky130_fd_sc_hd__conb_1 user_proj_example_71 (.LO(net71));
 sky130_fd_sc_hd__conb_1 user_proj_example_72 (.LO(net72));
 sky130_fd_sc_hd__conb_1 user_proj_example_73 (.LO(net73));
 sky130_fd_sc_hd__conb_1 user_proj_example_74 (.LO(net74));
 sky130_fd_sc_hd__conb_1 user_proj_example_75 (.LO(net75));
 sky130_fd_sc_hd__conb_1 user_proj_example_76 (.LO(net76));
 sky130_fd_sc_hd__conb_1 user_proj_example_77 (.LO(net77));
 sky130_fd_sc_hd__conb_1 user_proj_example_78 (.LO(net78));
 sky130_fd_sc_hd__conb_1 user_proj_example_79 (.LO(net79));
 sky130_fd_sc_hd__conb_1 user_proj_example_80 (.LO(net80));
 sky130_fd_sc_hd__conb_1 user_proj_example_81 (.LO(net81));
 sky130_fd_sc_hd__conb_1 user_proj_example_82 (.LO(net82));
 sky130_fd_sc_hd__conb_1 user_proj_example_83 (.LO(net83));
 sky130_fd_sc_hd__conb_1 user_proj_example_84 (.LO(net84));
 sky130_fd_sc_hd__conb_1 user_proj_example_85 (.LO(net85));
 sky130_fd_sc_hd__conb_1 user_proj_example_86 (.LO(net86));
 sky130_fd_sc_hd__conb_1 user_proj_example_87 (.LO(net87));
 sky130_fd_sc_hd__conb_1 user_proj_example_88 (.LO(net88));
 sky130_fd_sc_hd__conb_1 user_proj_example_89 (.LO(net89));
 sky130_fd_sc_hd__conb_1 user_proj_example_90 (.LO(net90));
 sky130_fd_sc_hd__conb_1 user_proj_example_91 (.LO(net91));
 sky130_fd_sc_hd__conb_1 user_proj_example_92 (.LO(net92));
 sky130_fd_sc_hd__conb_1 user_proj_example_93 (.LO(net93));
 sky130_fd_sc_hd__conb_1 user_proj_example_94 (.LO(net94));
 sky130_fd_sc_hd__conb_1 user_proj_example_95 (.LO(net95));
 sky130_fd_sc_hd__conb_1 user_proj_example_96 (.LO(net96));
 sky130_fd_sc_hd__conb_1 user_proj_example_97 (.LO(net97));
 sky130_fd_sc_hd__conb_1 user_proj_example_98 (.LO(net98));
 sky130_fd_sc_hd__conb_1 user_proj_example_99 (.LO(net99));
 sky130_fd_sc_hd__conb_1 user_proj_example_100 (.LO(net100));
 sky130_fd_sc_hd__conb_1 user_proj_example_101 (.LO(net101));
 sky130_fd_sc_hd__conb_1 user_proj_example_102 (.LO(net102));
 sky130_fd_sc_hd__conb_1 user_proj_example_103 (.LO(net103));
 sky130_fd_sc_hd__conb_1 user_proj_example_104 (.LO(net104));
 sky130_fd_sc_hd__conb_1 user_proj_example_105 (.LO(net105));
 sky130_fd_sc_hd__conb_1 user_proj_example_106 (.LO(net106));
 sky130_fd_sc_hd__conb_1 user_proj_example_107 (.LO(net107));
 sky130_fd_sc_hd__conb_1 user_proj_example_108 (.LO(net108));
 sky130_fd_sc_hd__conb_1 user_proj_example_109 (.LO(net109));
 sky130_fd_sc_hd__conb_1 user_proj_example_110 (.LO(net110));
 sky130_fd_sc_hd__conb_1 user_proj_example_111 (.LO(net111));
 sky130_fd_sc_hd__conb_1 user_proj_example_112 (.LO(net112));
 sky130_fd_sc_hd__conb_1 user_proj_example_113 (.LO(net113));
 sky130_fd_sc_hd__conb_1 user_proj_example_114 (.LO(net114));
 sky130_fd_sc_hd__conb_1 user_proj_example_115 (.LO(net115));
 sky130_fd_sc_hd__conb_1 user_proj_example_116 (.LO(net116));
 sky130_fd_sc_hd__conb_1 user_proj_example_117 (.LO(net117));
 sky130_fd_sc_hd__conb_1 user_proj_example_118 (.LO(net118));
 sky130_fd_sc_hd__conb_1 user_proj_example_119 (.LO(net119));
 sky130_fd_sc_hd__conb_1 user_proj_example_120 (.LO(net120));
 sky130_fd_sc_hd__conb_1 user_proj_example_121 (.LO(net121));
 sky130_fd_sc_hd__conb_1 user_proj_example_122 (.LO(net122));
 sky130_fd_sc_hd__conb_1 user_proj_example_123 (.LO(net123));
 sky130_fd_sc_hd__conb_1 user_proj_example_124 (.LO(net124));
 sky130_fd_sc_hd__conb_1 user_proj_example_125 (.LO(net125));
 sky130_fd_sc_hd__conb_1 user_proj_example_126 (.LO(net126));
 sky130_fd_sc_hd__conb_1 user_proj_example_127 (.LO(net127));
 sky130_fd_sc_hd__conb_1 user_proj_example_128 (.LO(net128));
 sky130_fd_sc_hd__conb_1 user_proj_example_129 (.LO(net129));
 sky130_fd_sc_hd__conb_1 user_proj_example_130 (.LO(net130));
 sky130_fd_sc_hd__conb_1 user_proj_example_131 (.LO(net131));
 sky130_fd_sc_hd__conb_1 user_proj_example_132 (.LO(net132));
 sky130_fd_sc_hd__conb_1 user_proj_example_133 (.LO(net133));
 sky130_fd_sc_hd__conb_1 user_proj_example_134 (.LO(net134));
 sky130_fd_sc_hd__conb_1 user_proj_example_135 (.LO(net135));
 sky130_fd_sc_hd__conb_1 user_proj_example_136 (.LO(net136));
 sky130_fd_sc_hd__conb_1 user_proj_example_137 (.LO(net137));
 sky130_fd_sc_hd__conb_1 user_proj_example_138 (.LO(net138));
 sky130_fd_sc_hd__conb_1 user_proj_example_139 (.LO(net139));
 sky130_fd_sc_hd__conb_1 user_proj_example_140 (.LO(net140));
 sky130_fd_sc_hd__conb_1 user_proj_example_141 (.LO(net141));
 sky130_fd_sc_hd__conb_1 user_proj_example_142 (.LO(net142));
 sky130_fd_sc_hd__conb_1 user_proj_example_143 (.LO(net143));
 sky130_fd_sc_hd__conb_1 user_proj_example_144 (.LO(net144));
 sky130_fd_sc_hd__conb_1 user_proj_example_145 (.LO(net145));
 sky130_fd_sc_hd__conb_1 user_proj_example_146 (.LO(net146));
 sky130_fd_sc_hd__conb_1 user_proj_example_147 (.LO(net147));
 sky130_fd_sc_hd__conb_1 user_proj_example_148 (.LO(net148));
 sky130_fd_sc_hd__conb_1 user_proj_example_149 (.LO(net149));
 sky130_fd_sc_hd__conb_1 user_proj_example_150 (.LO(net150));
 sky130_fd_sc_hd__conb_1 user_proj_example_151 (.LO(net151));
 sky130_fd_sc_hd__conb_1 user_proj_example_152 (.LO(net152));
 sky130_fd_sc_hd__conb_1 user_proj_example_153 (.LO(net153));
 sky130_fd_sc_hd__conb_1 user_proj_example_154 (.LO(net154));
 sky130_fd_sc_hd__conb_1 user_proj_example_155 (.LO(net155));
 sky130_fd_sc_hd__conb_1 user_proj_example_156 (.LO(net156));
 sky130_fd_sc_hd__conb_1 user_proj_example_157 (.LO(net157));
 sky130_fd_sc_hd__conb_1 user_proj_example_158 (.LO(net158));
 sky130_fd_sc_hd__conb_1 user_proj_example_159 (.LO(net159));
 sky130_fd_sc_hd__conb_1 user_proj_example_160 (.LO(net160));
 sky130_fd_sc_hd__conb_1 user_proj_example_161 (.LO(net161));
 sky130_fd_sc_hd__conb_1 user_proj_example_162 (.LO(net162));
 sky130_fd_sc_hd__conb_1 user_proj_example_163 (.LO(net163));
 sky130_fd_sc_hd__conb_1 user_proj_example_164 (.LO(net164));
 sky130_fd_sc_hd__conb_1 user_proj_example_165 (.LO(net165));
 sky130_fd_sc_hd__conb_1 user_proj_example_166 (.LO(net166));
 sky130_fd_sc_hd__conb_1 user_proj_example_167 (.LO(net167));
 sky130_fd_sc_hd__conb_1 user_proj_example_168 (.LO(net168));
 sky130_fd_sc_hd__conb_1 user_proj_example_169 (.LO(net169));
 sky130_fd_sc_hd__conb_1 user_proj_example_170 (.LO(net170));
 sky130_fd_sc_hd__conb_1 user_proj_example_171 (.LO(net171));
 sky130_fd_sc_hd__conb_1 user_proj_example_172 (.LO(net172));
 sky130_fd_sc_hd__conb_1 user_proj_example_173 (.LO(net173));
 sky130_fd_sc_hd__conb_1 user_proj_example_174 (.LO(net174));
 sky130_fd_sc_hd__conb_1 user_proj_example_175 (.LO(net175));
 sky130_fd_sc_hd__conb_1 user_proj_example_176 (.LO(net176));
 sky130_fd_sc_hd__conb_1 user_proj_example_177 (.LO(net177));
 sky130_fd_sc_hd__conb_1 user_proj_example_178 (.LO(net178));
 sky130_fd_sc_hd__conb_1 user_proj_example_179 (.LO(net179));
 sky130_fd_sc_hd__conb_1 user_proj_example_180 (.LO(net180));
 sky130_fd_sc_hd__conb_1 user_proj_example_181 (.LO(net181));
 sky130_fd_sc_hd__conb_1 user_proj_example_182 (.LO(net182));
 sky130_fd_sc_hd__conb_1 user_proj_example_183 (.LO(net183));
 sky130_fd_sc_hd__conb_1 user_proj_example_184 (.LO(net184));
 sky130_fd_sc_hd__conb_1 user_proj_example_185 (.LO(net185));
 sky130_fd_sc_hd__conb_1 user_proj_example_186 (.LO(net186));
 sky130_fd_sc_hd__conb_1 user_proj_example_187 (.LO(net187));
 sky130_fd_sc_hd__conb_1 user_proj_example_188 (.LO(net188));
 sky130_fd_sc_hd__conb_1 user_proj_example_189 (.LO(net189));
 sky130_fd_sc_hd__conb_1 user_proj_example_190 (.LO(net190));
 sky130_fd_sc_hd__conb_1 user_proj_example_191 (.LO(net191));
 sky130_fd_sc_hd__conb_1 user_proj_example_192 (.LO(net192));
 sky130_fd_sc_hd__conb_1 user_proj_example_193 (.LO(net193));
 sky130_fd_sc_hd__conb_1 user_proj_example_194 (.LO(net194));
 sky130_fd_sc_hd__conb_1 user_proj_example_195 (.LO(net195));
 sky130_fd_sc_hd__conb_1 user_proj_example_196 (.LO(net196));
 sky130_fd_sc_hd__conb_1 user_proj_example_197 (.LO(net197));
 sky130_fd_sc_hd__conb_1 user_proj_example_198 (.LO(net198));
 sky130_fd_sc_hd__conb_1 user_proj_example_199 (.LO(net199));
 sky130_fd_sc_hd__conb_1 user_proj_example_200 (.LO(net200));
 sky130_fd_sc_hd__conb_1 user_proj_example_201 (.LO(net201));
 sky130_fd_sc_hd__conb_1 user_proj_example_202 (.LO(net202));
 sky130_fd_sc_hd__conb_1 user_proj_example_203 (.LO(net203));
 sky130_fd_sc_hd__conb_1 user_proj_example_204 (.LO(net204));
 sky130_fd_sc_hd__conb_1 user_proj_example_205 (.LO(net205));
 sky130_fd_sc_hd__conb_1 user_proj_example_206 (.LO(net206));
 sky130_fd_sc_hd__conb_1 user_proj_example_207 (.LO(net207));
 sky130_fd_sc_hd__conb_1 user_proj_example_208 (.LO(net208));
 sky130_fd_sc_hd__conb_1 user_proj_example_209 (.LO(net209));
 sky130_fd_sc_hd__conb_1 user_proj_example_210 (.LO(net210));
 sky130_fd_sc_hd__conb_1 user_proj_example_211 (.LO(net211));
 sky130_fd_sc_hd__conb_1 user_proj_example_212 (.LO(net212));
 sky130_fd_sc_hd__conb_1 user_proj_example_213 (.LO(net213));
 sky130_fd_sc_hd__conb_1 user_proj_example_214 (.LO(net214));
 sky130_fd_sc_hd__conb_1 user_proj_example_215 (.LO(net215));
 sky130_fd_sc_hd__conb_1 user_proj_example_216 (.LO(net216));
 sky130_fd_sc_hd__conb_1 user_proj_example_217 (.LO(net217));
 sky130_fd_sc_hd__conb_1 user_proj_example_218 (.LO(net218));
 sky130_fd_sc_hd__conb_1 user_proj_example_219 (.LO(net219));
 sky130_fd_sc_hd__conb_1 user_proj_example_220 (.LO(net220));
 sky130_fd_sc_hd__conb_1 user_proj_example_221 (.LO(net221));
 sky130_fd_sc_hd__conb_1 user_proj_example_222 (.LO(net222));
 sky130_fd_sc_hd__conb_1 user_proj_example_223 (.LO(net223));
 sky130_fd_sc_hd__conb_1 user_proj_example_224 (.LO(net224));
 sky130_fd_sc_hd__conb_1 user_proj_example_225 (.LO(net225));
 sky130_fd_sc_hd__conb_1 user_proj_example_226 (.LO(net226));
 sky130_fd_sc_hd__conb_1 user_proj_example_227 (.LO(net227));
 sky130_fd_sc_hd__conb_1 user_proj_example_228 (.LO(net228));
 sky130_fd_sc_hd__conb_1 user_proj_example_229 (.LO(net229));
 sky130_fd_sc_hd__conb_1 user_proj_example_230 (.LO(net230));
 sky130_fd_sc_hd__conb_1 user_proj_example_231 (.LO(net231));
 sky130_fd_sc_hd__conb_1 user_proj_example_232 (.LO(net232));
 sky130_fd_sc_hd__conb_1 user_proj_example_233 (.LO(net233));
 sky130_fd_sc_hd__conb_1 user_proj_example_234 (.LO(net234));
 sky130_fd_sc_hd__conb_1 user_proj_example_235 (.LO(net235));
 sky130_fd_sc_hd__conb_1 user_proj_example_236 (.LO(net236));
 sky130_fd_sc_hd__conb_1 user_proj_example_237 (.LO(net237));
 sky130_fd_sc_hd__conb_1 user_proj_example_238 (.LO(net238));
 sky130_fd_sc_hd__conb_1 user_proj_example_239 (.LO(net239));
 sky130_fd_sc_hd__conb_1 user_proj_example_240 (.LO(net240));
 sky130_fd_sc_hd__conb_1 user_proj_example_241 (.LO(net241));
 sky130_fd_sc_hd__conb_1 user_proj_example_242 (.LO(net242));
 sky130_fd_sc_hd__conb_1 user_proj_example_243 (.LO(net243));
 sky130_fd_sc_hd__conb_1 user_proj_example_244 (.LO(net244));
 sky130_fd_sc_hd__conb_1 user_proj_example_245 (.LO(net245));
 sky130_fd_sc_hd__conb_1 user_proj_example_246 (.LO(net246));
 sky130_fd_sc_hd__conb_1 user_proj_example_247 (.LO(net247));
 sky130_fd_sc_hd__conb_1 user_proj_example_248 (.LO(net248));
 sky130_fd_sc_hd__conb_1 user_proj_example_249 (.LO(net249));
 sky130_fd_sc_hd__conb_1 user_proj_example_250 (.LO(net250));
 sky130_fd_sc_hd__conb_1 user_proj_example_251 (.LO(net251));
 sky130_fd_sc_hd__conb_1 user_proj_example_252 (.LO(net252));
 sky130_fd_sc_hd__conb_1 user_proj_example_253 (.LO(net253));
 sky130_fd_sc_hd__conb_1 user_proj_example_254 (.LO(net254));
 sky130_fd_sc_hd__conb_1 user_proj_example_255 (.LO(net255));
 sky130_fd_sc_hd__conb_1 user_proj_example_256 (.LO(net256));
 sky130_fd_sc_hd__conb_1 user_proj_example_257 (.LO(net257));
 sky130_fd_sc_hd__conb_1 user_proj_example_258 (.LO(net258));
 sky130_fd_sc_hd__conb_1 user_proj_example_259 (.LO(net259));
 sky130_fd_sc_hd__conb_1 user_proj_example_260 (.LO(net260));
 sky130_fd_sc_hd__conb_1 user_proj_example_261 (.LO(net261));
 sky130_fd_sc_hd__conb_1 user_proj_example_262 (.LO(net262));
 sky130_fd_sc_hd__conb_1 _4237__263 (.HI(net263));
 sky130_fd_sc_hd__clkbuf_1 _4873_ (.A(net6),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_1 _4874_ (.A(net1),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_1 _4875_ (.A(net2),
    .X(net9));
 sky130_fd_sc_hd__ebufn_2 _4876_ (.A(\usb2uart.dn_tx ),
    .TE_B(_2085_),
    .Z(net1));
 sky130_fd_sc_hd__ebufn_2 _4877_ (.A(\usb2uart.dp_tx ),
    .TE_B(_2086_),
    .Z(net2));
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__decap_3 PHY_130 ();
 sky130_fd_sc_hd__decap_3 PHY_131 ();
 sky130_fd_sc_hd__decap_3 PHY_132 ();
 sky130_fd_sc_hd__decap_3 PHY_133 ();
 sky130_fd_sc_hd__decap_3 PHY_134 ();
 sky130_fd_sc_hd__decap_3 PHY_135 ();
 sky130_fd_sc_hd__decap_3 PHY_136 ();
 sky130_fd_sc_hd__decap_3 PHY_137 ();
 sky130_fd_sc_hd__decap_3 PHY_138 ();
 sky130_fd_sc_hd__decap_3 PHY_139 ();
 sky130_fd_sc_hd__decap_3 PHY_140 ();
 sky130_fd_sc_hd__decap_3 PHY_141 ();
 sky130_fd_sc_hd__decap_3 PHY_142 ();
 sky130_fd_sc_hd__decap_3 PHY_143 ();
 sky130_fd_sc_hd__decap_3 PHY_144 ();
 sky130_fd_sc_hd__decap_3 PHY_145 ();
 sky130_fd_sc_hd__decap_3 PHY_146 ();
 sky130_fd_sc_hd__decap_3 PHY_147 ();
 sky130_fd_sc_hd__decap_3 PHY_148 ();
 sky130_fd_sc_hd__decap_3 PHY_149 ();
 sky130_fd_sc_hd__decap_3 PHY_150 ();
 sky130_fd_sc_hd__decap_3 PHY_151 ();
 sky130_fd_sc_hd__decap_3 PHY_152 ();
 sky130_fd_sc_hd__decap_3 PHY_153 ();
 sky130_fd_sc_hd__decap_3 PHY_154 ();
 sky130_fd_sc_hd__decap_3 PHY_155 ();
 sky130_fd_sc_hd__decap_3 PHY_156 ();
 sky130_fd_sc_hd__decap_3 PHY_157 ();
 sky130_fd_sc_hd__decap_3 PHY_158 ();
 sky130_fd_sc_hd__decap_3 PHY_159 ();
 sky130_fd_sc_hd__decap_3 PHY_160 ();
 sky130_fd_sc_hd__decap_3 PHY_161 ();
 sky130_fd_sc_hd__decap_3 PHY_162 ();
 sky130_fd_sc_hd__decap_3 PHY_163 ();
 sky130_fd_sc_hd__decap_3 PHY_164 ();
 sky130_fd_sc_hd__decap_3 PHY_165 ();
 sky130_fd_sc_hd__decap_3 PHY_166 ();
 sky130_fd_sc_hd__decap_3 PHY_167 ();
 sky130_fd_sc_hd__decap_3 PHY_168 ();
 sky130_fd_sc_hd__decap_3 PHY_169 ();
 sky130_fd_sc_hd__decap_3 PHY_170 ();
 sky130_fd_sc_hd__decap_3 PHY_171 ();
 sky130_fd_sc_hd__decap_3 PHY_172 ();
 sky130_fd_sc_hd__decap_3 PHY_173 ();
 sky130_fd_sc_hd__decap_3 PHY_174 ();
 sky130_fd_sc_hd__decap_3 PHY_175 ();
 sky130_fd_sc_hd__decap_3 PHY_176 ();
 sky130_fd_sc_hd__decap_3 PHY_177 ();
 sky130_fd_sc_hd__decap_3 PHY_178 ();
 sky130_fd_sc_hd__decap_3 PHY_179 ();
 sky130_fd_sc_hd__decap_3 PHY_180 ();
 sky130_fd_sc_hd__decap_3 PHY_181 ();
 sky130_fd_sc_hd__decap_3 PHY_182 ();
 sky130_fd_sc_hd__decap_3 PHY_183 ();
 sky130_fd_sc_hd__decap_3 PHY_184 ();
 sky130_fd_sc_hd__decap_3 PHY_185 ();
 sky130_fd_sc_hd__decap_3 PHY_186 ();
 sky130_fd_sc_hd__decap_3 PHY_187 ();
 sky130_fd_sc_hd__decap_3 PHY_188 ();
 sky130_fd_sc_hd__decap_3 PHY_189 ();
 sky130_fd_sc_hd__decap_3 PHY_190 ();
 sky130_fd_sc_hd__decap_3 PHY_191 ();
 sky130_fd_sc_hd__decap_3 PHY_192 ();
 sky130_fd_sc_hd__decap_3 PHY_193 ();
 sky130_fd_sc_hd__decap_3 PHY_194 ();
 sky130_fd_sc_hd__decap_3 PHY_195 ();
 sky130_fd_sc_hd__decap_3 PHY_196 ();
 sky130_fd_sc_hd__decap_3 PHY_197 ();
 sky130_fd_sc_hd__decap_3 PHY_198 ();
 sky130_fd_sc_hd__decap_3 PHY_199 ();
 sky130_fd_sc_hd__decap_3 PHY_200 ();
 sky130_fd_sc_hd__decap_3 PHY_201 ();
 sky130_fd_sc_hd__decap_3 PHY_202 ();
 sky130_fd_sc_hd__decap_3 PHY_203 ();
 sky130_fd_sc_hd__decap_3 PHY_204 ();
 sky130_fd_sc_hd__decap_3 PHY_205 ();
 sky130_fd_sc_hd__decap_3 PHY_206 ();
 sky130_fd_sc_hd__decap_3 PHY_207 ();
 sky130_fd_sc_hd__decap_3 PHY_208 ();
 sky130_fd_sc_hd__decap_3 PHY_209 ();
 sky130_fd_sc_hd__decap_3 PHY_210 ();
 sky130_fd_sc_hd__decap_3 PHY_211 ();
 sky130_fd_sc_hd__decap_3 PHY_212 ();
 sky130_fd_sc_hd__decap_3 PHY_213 ();
 sky130_fd_sc_hd__decap_3 PHY_214 ();
 sky130_fd_sc_hd__decap_3 PHY_215 ();
 sky130_fd_sc_hd__decap_3 PHY_216 ();
 sky130_fd_sc_hd__decap_3 PHY_217 ();
 sky130_fd_sc_hd__decap_3 PHY_218 ();
 sky130_fd_sc_hd__decap_3 PHY_219 ();
 sky130_fd_sc_hd__decap_3 PHY_220 ();
 sky130_fd_sc_hd__decap_3 PHY_221 ();
 sky130_fd_sc_hd__decap_3 PHY_222 ();
 sky130_fd_sc_hd__decap_3 PHY_223 ();
 sky130_fd_sc_hd__decap_3 PHY_224 ();
 sky130_fd_sc_hd__decap_3 PHY_225 ();
 sky130_fd_sc_hd__decap_3 PHY_226 ();
 sky130_fd_sc_hd__decap_3 PHY_227 ();
 sky130_fd_sc_hd__decap_3 PHY_228 ();
 sky130_fd_sc_hd__decap_3 PHY_229 ();
 sky130_fd_sc_hd__decap_3 PHY_230 ();
 sky130_fd_sc_hd__decap_3 PHY_231 ();
 sky130_fd_sc_hd__decap_3 PHY_232 ();
 sky130_fd_sc_hd__decap_3 PHY_233 ();
 sky130_fd_sc_hd__decap_3 PHY_234 ();
 sky130_fd_sc_hd__decap_3 PHY_235 ();
 sky130_fd_sc_hd__decap_3 PHY_236 ();
 sky130_fd_sc_hd__decap_3 PHY_237 ();
 sky130_fd_sc_hd__decap_3 PHY_238 ();
 sky130_fd_sc_hd__decap_3 PHY_239 ();
 sky130_fd_sc_hd__decap_3 PHY_240 ();
 sky130_fd_sc_hd__decap_3 PHY_241 ();
 sky130_fd_sc_hd__decap_3 PHY_242 ();
 sky130_fd_sc_hd__decap_3 PHY_243 ();
 sky130_fd_sc_hd__decap_3 PHY_244 ();
 sky130_fd_sc_hd__decap_3 PHY_245 ();
 sky130_fd_sc_hd__decap_3 PHY_246 ();
 sky130_fd_sc_hd__decap_3 PHY_247 ();
 sky130_fd_sc_hd__decap_3 PHY_248 ();
 sky130_fd_sc_hd__decap_3 PHY_249 ();
 sky130_fd_sc_hd__decap_3 PHY_250 ();
 sky130_fd_sc_hd__decap_3 PHY_251 ();
 sky130_fd_sc_hd__decap_3 PHY_252 ();
 sky130_fd_sc_hd__decap_3 PHY_253 ();
 sky130_fd_sc_hd__decap_3 PHY_254 ();
 sky130_fd_sc_hd__decap_3 PHY_255 ();
 sky130_fd_sc_hd__decap_3 PHY_256 ();
 sky130_fd_sc_hd__decap_3 PHY_257 ();
 sky130_fd_sc_hd__decap_3 PHY_258 ();
 sky130_fd_sc_hd__decap_3 PHY_259 ();
 sky130_fd_sc_hd__decap_3 PHY_260 ();
 sky130_fd_sc_hd__decap_3 PHY_261 ();
 sky130_fd_sc_hd__decap_3 PHY_262 ();
 sky130_fd_sc_hd__decap_3 PHY_263 ();
 sky130_fd_sc_hd__decap_3 PHY_264 ();
 sky130_fd_sc_hd__decap_3 PHY_265 ();
 sky130_fd_sc_hd__decap_3 PHY_266 ();
 sky130_fd_sc_hd__decap_3 PHY_267 ();
 sky130_fd_sc_hd__decap_3 PHY_268 ();
 sky130_fd_sc_hd__decap_3 PHY_269 ();
 sky130_fd_sc_hd__decap_3 PHY_270 ();
 sky130_fd_sc_hd__decap_3 PHY_271 ();
 sky130_fd_sc_hd__decap_3 PHY_272 ();
 sky130_fd_sc_hd__decap_3 PHY_273 ();
 sky130_fd_sc_hd__decap_3 PHY_274 ();
 sky130_fd_sc_hd__decap_3 PHY_275 ();
 sky130_fd_sc_hd__decap_3 PHY_276 ();
 sky130_fd_sc_hd__decap_3 PHY_277 ();
 sky130_fd_sc_hd__decap_3 PHY_278 ();
 sky130_fd_sc_hd__decap_3 PHY_279 ();
 sky130_fd_sc_hd__decap_3 PHY_280 ();
 sky130_fd_sc_hd__decap_3 PHY_281 ();
 sky130_fd_sc_hd__decap_3 PHY_282 ();
 sky130_fd_sc_hd__decap_3 PHY_283 ();
 sky130_fd_sc_hd__decap_3 PHY_284 ();
 sky130_fd_sc_hd__decap_3 PHY_285 ();
 sky130_fd_sc_hd__decap_3 PHY_286 ();
 sky130_fd_sc_hd__decap_3 PHY_287 ();
 sky130_fd_sc_hd__decap_3 PHY_288 ();
 sky130_fd_sc_hd__decap_3 PHY_289 ();
 sky130_fd_sc_hd__decap_3 PHY_290 ();
 sky130_fd_sc_hd__decap_3 PHY_291 ();
 sky130_fd_sc_hd__decap_3 PHY_292 ();
 sky130_fd_sc_hd__decap_3 PHY_293 ();
 sky130_fd_sc_hd__decap_3 PHY_294 ();
 sky130_fd_sc_hd__decap_3 PHY_295 ();
 sky130_fd_sc_hd__decap_3 PHY_296 ();
 sky130_fd_sc_hd__decap_3 PHY_297 ();
 sky130_fd_sc_hd__decap_3 PHY_298 ();
 sky130_fd_sc_hd__decap_3 PHY_299 ();
 sky130_fd_sc_hd__decap_3 PHY_300 ();
 sky130_fd_sc_hd__decap_3 PHY_301 ();
 sky130_fd_sc_hd__decap_3 PHY_302 ();
 sky130_fd_sc_hd__decap_3 PHY_303 ();
 sky130_fd_sc_hd__decap_3 PHY_304 ();
 sky130_fd_sc_hd__decap_3 PHY_305 ();
 sky130_fd_sc_hd__decap_3 PHY_306 ();
 sky130_fd_sc_hd__decap_3 PHY_307 ();
 sky130_fd_sc_hd__decap_3 PHY_308 ();
 sky130_fd_sc_hd__decap_3 PHY_309 ();
 sky130_fd_sc_hd__decap_3 PHY_310 ();
 sky130_fd_sc_hd__decap_3 PHY_311 ();
 sky130_fd_sc_hd__decap_3 PHY_312 ();
 sky130_fd_sc_hd__decap_3 PHY_313 ();
 sky130_fd_sc_hd__decap_3 PHY_314 ();
 sky130_fd_sc_hd__decap_3 PHY_315 ();
 sky130_fd_sc_hd__decap_3 PHY_316 ();
 sky130_fd_sc_hd__decap_3 PHY_317 ();
 sky130_fd_sc_hd__decap_3 PHY_318 ();
 sky130_fd_sc_hd__decap_3 PHY_319 ();
 sky130_fd_sc_hd__decap_3 PHY_320 ();
 sky130_fd_sc_hd__decap_3 PHY_321 ();
 sky130_fd_sc_hd__decap_3 PHY_322 ();
 sky130_fd_sc_hd__decap_3 PHY_323 ();
 sky130_fd_sc_hd__decap_3 PHY_324 ();
 sky130_fd_sc_hd__decap_3 PHY_325 ();
 sky130_fd_sc_hd__decap_3 PHY_326 ();
 sky130_fd_sc_hd__decap_3 PHY_327 ();
 sky130_fd_sc_hd__decap_3 PHY_328 ();
 sky130_fd_sc_hd__decap_3 PHY_329 ();
 sky130_fd_sc_hd__decap_3 PHY_330 ();
 sky130_fd_sc_hd__decap_3 PHY_331 ();
 sky130_fd_sc_hd__decap_3 PHY_332 ();
 sky130_fd_sc_hd__decap_3 PHY_333 ();
 sky130_fd_sc_hd__decap_3 PHY_334 ();
 sky130_fd_sc_hd__decap_3 PHY_335 ();
 sky130_fd_sc_hd__decap_3 PHY_336 ();
 sky130_fd_sc_hd__decap_3 PHY_337 ();
 sky130_fd_sc_hd__decap_3 PHY_338 ();
 sky130_fd_sc_hd__decap_3 PHY_339 ();
 sky130_fd_sc_hd__decap_3 PHY_340 ();
 sky130_fd_sc_hd__decap_3 PHY_341 ();
 sky130_fd_sc_hd__decap_3 PHY_342 ();
 sky130_fd_sc_hd__decap_3 PHY_343 ();
 sky130_fd_sc_hd__decap_3 PHY_344 ();
 sky130_fd_sc_hd__decap_3 PHY_345 ();
 sky130_fd_sc_hd__decap_3 PHY_346 ();
 sky130_fd_sc_hd__decap_3 PHY_347 ();
 sky130_fd_sc_hd__decap_3 PHY_348 ();
 sky130_fd_sc_hd__decap_3 PHY_349 ();
 sky130_fd_sc_hd__decap_3 PHY_350 ();
 sky130_fd_sc_hd__decap_3 PHY_351 ();
 sky130_fd_sc_hd__decap_3 PHY_352 ();
 sky130_fd_sc_hd__decap_3 PHY_353 ();
 sky130_fd_sc_hd__decap_3 PHY_354 ();
 sky130_fd_sc_hd__decap_3 PHY_355 ();
 sky130_fd_sc_hd__decap_3 PHY_356 ();
 sky130_fd_sc_hd__decap_3 PHY_357 ();
 sky130_fd_sc_hd__decap_3 PHY_358 ();
 sky130_fd_sc_hd__decap_3 PHY_359 ();
 sky130_fd_sc_hd__decap_3 PHY_360 ();
 sky130_fd_sc_hd__decap_3 PHY_361 ();
 sky130_fd_sc_hd__decap_3 PHY_362 ();
 sky130_fd_sc_hd__decap_3 PHY_363 ();
 sky130_fd_sc_hd__decap_3 PHY_364 ();
 sky130_fd_sc_hd__decap_3 PHY_365 ();
 sky130_fd_sc_hd__decap_3 PHY_366 ();
 sky130_fd_sc_hd__decap_3 PHY_367 ();
 sky130_fd_sc_hd__decap_3 PHY_368 ();
 sky130_fd_sc_hd__decap_3 PHY_369 ();
 sky130_fd_sc_hd__decap_3 PHY_370 ();
 sky130_fd_sc_hd__decap_3 PHY_371 ();
 sky130_fd_sc_hd__decap_3 PHY_372 ();
 sky130_fd_sc_hd__decap_3 PHY_373 ();
 sky130_fd_sc_hd__decap_3 PHY_374 ();
 sky130_fd_sc_hd__decap_3 PHY_375 ();
 sky130_fd_sc_hd__decap_3 PHY_376 ();
 sky130_fd_sc_hd__decap_3 PHY_377 ();
 sky130_fd_sc_hd__decap_3 PHY_378 ();
 sky130_fd_sc_hd__decap_3 PHY_379 ();
 sky130_fd_sc_hd__decap_3 PHY_380 ();
 sky130_fd_sc_hd__decap_3 PHY_381 ();
 sky130_fd_sc_hd__decap_3 PHY_382 ();
 sky130_fd_sc_hd__decap_3 PHY_383 ();
 sky130_fd_sc_hd__decap_3 PHY_384 ();
 sky130_fd_sc_hd__decap_3 PHY_385 ();
 sky130_fd_sc_hd__decap_3 PHY_386 ();
 sky130_fd_sc_hd__decap_3 PHY_387 ();
 sky130_fd_sc_hd__decap_3 PHY_388 ();
 sky130_fd_sc_hd__decap_3 PHY_389 ();
 sky130_fd_sc_hd__decap_3 PHY_390 ();
 sky130_fd_sc_hd__decap_3 PHY_391 ();
 sky130_fd_sc_hd__decap_3 PHY_392 ();
 sky130_fd_sc_hd__decap_3 PHY_393 ();
 sky130_fd_sc_hd__decap_3 PHY_394 ();
 sky130_fd_sc_hd__decap_3 PHY_395 ();
 sky130_fd_sc_hd__decap_3 PHY_396 ();
 sky130_fd_sc_hd__decap_3 PHY_397 ();
 sky130_fd_sc_hd__decap_3 PHY_398 ();
 sky130_fd_sc_hd__decap_3 PHY_399 ();
 sky130_fd_sc_hd__decap_3 PHY_400 ();
 sky130_fd_sc_hd__decap_3 PHY_401 ();
 sky130_fd_sc_hd__decap_3 PHY_402 ();
 sky130_fd_sc_hd__decap_3 PHY_403 ();
 sky130_fd_sc_hd__decap_3 PHY_404 ();
 sky130_fd_sc_hd__decap_3 PHY_405 ();
 sky130_fd_sc_hd__decap_3 PHY_406 ();
 sky130_fd_sc_hd__decap_3 PHY_407 ();
 sky130_fd_sc_hd__decap_3 PHY_408 ();
 sky130_fd_sc_hd__decap_3 PHY_409 ();
 sky130_fd_sc_hd__decap_3 PHY_410 ();
 sky130_fd_sc_hd__decap_3 PHY_411 ();
 sky130_fd_sc_hd__decap_3 PHY_412 ();
 sky130_fd_sc_hd__decap_3 PHY_413 ();
 sky130_fd_sc_hd__decap_3 PHY_414 ();
 sky130_fd_sc_hd__decap_3 PHY_415 ();
 sky130_fd_sc_hd__decap_3 PHY_416 ();
 sky130_fd_sc_hd__decap_3 PHY_417 ();
 sky130_fd_sc_hd__decap_3 PHY_418 ();
 sky130_fd_sc_hd__decap_3 PHY_419 ();
 sky130_fd_sc_hd__decap_3 PHY_420 ();
 sky130_fd_sc_hd__decap_3 PHY_421 ();
 sky130_fd_sc_hd__decap_3 PHY_422 ();
 sky130_fd_sc_hd__decap_3 PHY_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7699 ();
 sky130_fd_sc_hd__clkbuf_2 input1 (.A(io_in[17]),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_2 input2 (.A(io_in[18]),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_2 input3 (.A(io_in[19]),
    .X(net3));
 sky130_fd_sc_hd__buf_8 input4 (.A(wb_rst_i),
    .X(net4));
 sky130_fd_sc_hd__buf_2 output5 (.A(net5),
    .X(io_oeb[17]));
 sky130_fd_sc_hd__buf_2 output6 (.A(net6),
    .X(io_oeb[18]));
 sky130_fd_sc_hd__buf_2 output7 (.A(net7),
    .X(io_out[16]));
 sky130_fd_sc_hd__buf_2 output8 (.A(net8),
    .X(io_out[17]));
 sky130_fd_sc_hd__buf_2 output9 (.A(net9),
    .X(io_out[18]));
 sky130_fd_sc_hd__buf_2 output10 (.A(net10),
    .X(io_out[20]));
 sky130_fd_sc_hd__clkbuf_4 fanout11 (.A(net12),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_4 fanout12 (.A(net15),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_4 fanout13 (.A(net15),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_2 fanout14 (.A(net15),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_2 fanout15 (.A(net22),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_4 fanout16 (.A(net18),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_4 fanout17 (.A(net18),
    .X(net17));
 sky130_fd_sc_hd__buf_2 fanout18 (.A(net22),
    .X(net18));
 sky130_fd_sc_hd__clkbuf_4 fanout19 (.A(net22),
    .X(net19));
 sky130_fd_sc_hd__buf_2 fanout20 (.A(net22),
    .X(net20));
 sky130_fd_sc_hd__clkbuf_4 fanout21 (.A(net22),
    .X(net21));
 sky130_fd_sc_hd__clkbuf_2 fanout22 (.A(net54),
    .X(net22));
 sky130_fd_sc_hd__clkbuf_4 fanout23 (.A(net25),
    .X(net23));
 sky130_fd_sc_hd__clkbuf_4 fanout24 (.A(net25),
    .X(net24));
 sky130_fd_sc_hd__buf_2 fanout25 (.A(net32),
    .X(net25));
 sky130_fd_sc_hd__clkbuf_4 fanout26 (.A(net32),
    .X(net26));
 sky130_fd_sc_hd__clkbuf_4 fanout27 (.A(net32),
    .X(net27));
 sky130_fd_sc_hd__clkbuf_4 fanout28 (.A(net30),
    .X(net28));
 sky130_fd_sc_hd__clkbuf_2 fanout29 (.A(net30),
    .X(net29));
 sky130_fd_sc_hd__clkbuf_2 fanout30 (.A(net32),
    .X(net30));
 sky130_fd_sc_hd__clkbuf_4 fanout31 (.A(net32),
    .X(net31));
 sky130_fd_sc_hd__buf_2 fanout32 (.A(net54),
    .X(net32));
 sky130_fd_sc_hd__clkbuf_4 fanout33 (.A(net34),
    .X(net33));
 sky130_fd_sc_hd__clkbuf_4 fanout34 (.A(net54),
    .X(net34));
 sky130_fd_sc_hd__clkbuf_4 fanout35 (.A(net38),
    .X(net35));
 sky130_fd_sc_hd__buf_2 fanout36 (.A(net38),
    .X(net36));
 sky130_fd_sc_hd__clkbuf_4 fanout37 (.A(net38),
    .X(net37));
 sky130_fd_sc_hd__clkbuf_2 fanout38 (.A(net54),
    .X(net38));
 sky130_fd_sc_hd__buf_4 fanout39 (.A(net43),
    .X(net39));
 sky130_fd_sc_hd__clkbuf_4 fanout40 (.A(net42),
    .X(net40));
 sky130_fd_sc_hd__clkbuf_4 fanout41 (.A(net43),
    .X(net41));
 sky130_fd_sc_hd__clkbuf_2 fanout42 (.A(net43),
    .X(net42));
 sky130_fd_sc_hd__buf_2 fanout43 (.A(net54),
    .X(net43));
 sky130_fd_sc_hd__clkbuf_4 fanout44 (.A(net46),
    .X(net44));
 sky130_fd_sc_hd__clkbuf_4 fanout45 (.A(net46),
    .X(net45));
 sky130_fd_sc_hd__clkbuf_4 fanout46 (.A(net53),
    .X(net46));
 sky130_fd_sc_hd__clkbuf_4 fanout47 (.A(net49),
    .X(net47));
 sky130_fd_sc_hd__buf_2 fanout48 (.A(net49),
    .X(net48));
 sky130_fd_sc_hd__clkbuf_4 fanout49 (.A(net53),
    .X(net49));
 sky130_fd_sc_hd__clkbuf_4 fanout50 (.A(net51),
    .X(net50));
 sky130_fd_sc_hd__buf_4 fanout51 (.A(net52),
    .X(net51));
 sky130_fd_sc_hd__clkbuf_4 fanout52 (.A(net53),
    .X(net52));
 sky130_fd_sc_hd__buf_2 fanout53 (.A(net54),
    .X(net53));
 sky130_fd_sc_hd__buf_4 fanout54 (.A(\usb2uart.u_usb_cdc.u_bulk_endp.rstn ),
    .X(net54));
 sky130_fd_sc_hd__clkbuf_4 fanout55 (.A(net56),
    .X(net55));
 sky130_fd_sc_hd__clkbuf_2 fanout56 (.A(net58),
    .X(net56));
 sky130_fd_sc_hd__clkbuf_4 fanout57 (.A(net58),
    .X(net57));
 sky130_fd_sc_hd__clkbuf_2 fanout58 (.A(net62),
    .X(net58));
 sky130_fd_sc_hd__clkbuf_4 fanout59 (.A(net61),
    .X(net59));
 sky130_fd_sc_hd__clkbuf_4 fanout60 (.A(net61),
    .X(net60));
 sky130_fd_sc_hd__buf_2 fanout61 (.A(net62),
    .X(net61));
 sky130_fd_sc_hd__buf_2 fanout62 (.A(net298),
    .X(net62));
 sky130_fd_sc_hd__conb_1 user_proj_example_63 (.LO(net63));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_1_user_clock2 (.A(clknet_2_0__leaf_user_clock2),
    .X(clknet_leaf_1_user_clock2));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_2_user_clock2 (.A(clknet_2_0__leaf_user_clock2),
    .X(clknet_leaf_2_user_clock2));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_3_user_clock2 (.A(clknet_2_0__leaf_user_clock2),
    .X(clknet_leaf_3_user_clock2));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_4_user_clock2 (.A(clknet_2_1__leaf_user_clock2),
    .X(clknet_leaf_4_user_clock2));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_5_user_clock2 (.A(clknet_2_0__leaf_user_clock2),
    .X(clknet_leaf_5_user_clock2));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_6_user_clock2 (.A(clknet_2_1__leaf_user_clock2),
    .X(clknet_leaf_6_user_clock2));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_8_user_clock2 (.A(clknet_2_1__leaf_user_clock2),
    .X(clknet_leaf_8_user_clock2));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_9_user_clock2 (.A(clknet_2_1__leaf_user_clock2),
    .X(clknet_leaf_9_user_clock2));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_10_user_clock2 (.A(clknet_2_1__leaf_user_clock2),
    .X(clknet_leaf_10_user_clock2));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_11_user_clock2 (.A(clknet_2_1__leaf_user_clock2),
    .X(clknet_leaf_11_user_clock2));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_12_user_clock2 (.A(clknet_2_1__leaf_user_clock2),
    .X(clknet_leaf_12_user_clock2));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_13_user_clock2 (.A(clknet_2_1__leaf_user_clock2),
    .X(clknet_leaf_13_user_clock2));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_14_user_clock2 (.A(clknet_2_3__leaf_user_clock2),
    .X(clknet_leaf_14_user_clock2));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_15_user_clock2 (.A(clknet_2_3__leaf_user_clock2),
    .X(clknet_leaf_15_user_clock2));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_16_user_clock2 (.A(clknet_2_3__leaf_user_clock2),
    .X(clknet_leaf_16_user_clock2));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_17_user_clock2 (.A(clknet_2_3__leaf_user_clock2),
    .X(clknet_leaf_17_user_clock2));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_18_user_clock2 (.A(clknet_2_3__leaf_user_clock2),
    .X(clknet_leaf_18_user_clock2));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_19_user_clock2 (.A(clknet_2_3__leaf_user_clock2),
    .X(clknet_leaf_19_user_clock2));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_20_user_clock2 (.A(clknet_2_3__leaf_user_clock2),
    .X(clknet_leaf_20_user_clock2));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_21_user_clock2 (.A(clknet_2_3__leaf_user_clock2),
    .X(clknet_leaf_21_user_clock2));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_22_user_clock2 (.A(clknet_2_2__leaf_user_clock2),
    .X(clknet_leaf_22_user_clock2));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_23_user_clock2 (.A(clknet_2_2__leaf_user_clock2),
    .X(clknet_leaf_23_user_clock2));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_24_user_clock2 (.A(clknet_opt_1_0_user_clock2),
    .X(clknet_leaf_24_user_clock2));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_25_user_clock2 (.A(clknet_2_2__leaf_user_clock2),
    .X(clknet_leaf_25_user_clock2));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_26_user_clock2 (.A(clknet_2_2__leaf_user_clock2),
    .X(clknet_leaf_26_user_clock2));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_27_user_clock2 (.A(clknet_2_2__leaf_user_clock2),
    .X(clknet_leaf_27_user_clock2));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_28_user_clock2 (.A(clknet_2_2__leaf_user_clock2),
    .X(clknet_leaf_28_user_clock2));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_29_user_clock2 (.A(clknet_2_2__leaf_user_clock2),
    .X(clknet_leaf_29_user_clock2));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_30_user_clock2 (.A(clknet_2_2__leaf_user_clock2),
    .X(clknet_leaf_30_user_clock2));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_31_user_clock2 (.A(clknet_2_2__leaf_user_clock2),
    .X(clknet_leaf_31_user_clock2));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_32_user_clock2 (.A(clknet_2_2__leaf_user_clock2),
    .X(clknet_leaf_32_user_clock2));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_33_user_clock2 (.A(clknet_2_0__leaf_user_clock2),
    .X(clknet_leaf_33_user_clock2));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_34_user_clock2 (.A(clknet_2_0__leaf_user_clock2),
    .X(clknet_leaf_34_user_clock2));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_35_user_clock2 (.A(clknet_2_0__leaf_user_clock2),
    .X(clknet_leaf_35_user_clock2));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_36_user_clock2 (.A(clknet_2_0__leaf_user_clock2),
    .X(clknet_leaf_36_user_clock2));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_37_user_clock2 (.A(clknet_2_0__leaf_user_clock2),
    .X(clknet_leaf_37_user_clock2));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_user_clock2 (.A(user_clock2),
    .X(clknet_0_user_clock2));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_0__f_user_clock2 (.A(clknet_0_user_clock2),
    .X(clknet_2_0__leaf_user_clock2));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_1__f_user_clock2 (.A(clknet_0_user_clock2),
    .X(clknet_2_1__leaf_user_clock2));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_2__f_user_clock2 (.A(clknet_0_user_clock2),
    .X(clknet_2_2__leaf_user_clock2));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_3__f_user_clock2 (.A(clknet_0_user_clock2),
    .X(clknet_2_3__leaf_user_clock2));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_opt_1_0_user_clock2 (.A(clknet_2_2__leaf_user_clock2),
    .X(clknet_opt_1_0_user_clock2));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1 (.A(\usb2uart.u_usb_cdc.rstn ),
    .X(net298));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2 (.A(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.dp_q[2] ),
    .X(net299));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3 (.A(\usb2uart.u_usb_cdc.u_sie.u_phy_rx.dn_q[2] ),
    .X(net300));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4 (.A(\usb2uart.u_usb_cdc.rstn_sq[1] ),
    .X(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA__4236__RESET_B (.DIODE(_0044_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4104__C1 (.DIODE(_0044_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4102__C1 (.DIODE(_0044_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4100__C1 (.DIODE(_0044_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4098__C1 (.DIODE(_0044_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4096__C1 (.DIODE(_0044_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4094__C1 (.DIODE(_0044_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4092__C1 (.DIODE(_0044_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4055__C1 (.DIODE(_0044_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4048__C1 (.DIODE(_0044_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3133__A (.DIODE(_0452_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3130__A_N (.DIODE(_0452_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3092__A2 (.DIODE(_0452_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3090__A (.DIODE(_0452_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3081__A (.DIODE(_0452_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3077__A (.DIODE(_0452_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3075__A (.DIODE(_0452_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2370__A (.DIODE(_0452_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2216__A (.DIODE(_0452_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2180__A (.DIODE(_0452_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3359__A1 (.DIODE(_0461_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2489__A1 (.DIODE(_0461_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2462__A1 (.DIODE(_0461_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2451__C (.DIODE(_0461_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2395__A1 (.DIODE(_0461_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2394__A1 (.DIODE(_0461_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2385__A1 (.DIODE(_0461_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2384__A (.DIODE(_0461_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2377__A (.DIODE(_0461_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2186__A (.DIODE(_0461_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3586__A1 (.DIODE(_0466_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3554__A (.DIODE(_0466_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3498__A1 (.DIODE(_0466_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2984__A (.DIODE(_0466_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2443__A_N (.DIODE(_0466_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2440__C1 (.DIODE(_0466_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2303__A (.DIODE(_0466_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2293__B (.DIODE(_0466_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2290__B (.DIODE(_0466_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2190__C (.DIODE(_0466_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3363__B1 (.DIODE(_0473_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3295__A1 (.DIODE(_0473_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3062__B1 (.DIODE(_0473_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2610__A1 (.DIODE(_0473_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2467__A1 (.DIODE(_0473_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2466__C1 (.DIODE(_0473_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2441__A (.DIODE(_0473_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2418__A (.DIODE(_0473_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2398__A2 (.DIODE(_0473_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2197__A (.DIODE(_0473_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3165__A1 (.DIODE(_0477_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3140__A1 (.DIODE(_0477_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3135__A2 (.DIODE(_0477_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2492__A (.DIODE(_0477_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2203__B (.DIODE(_0477_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2201__B (.DIODE(_0477_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3574__A1 (.DIODE(_0482_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3459__A (.DIODE(_0482_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2963__A (.DIODE(_0482_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2446__A (.DIODE(_0482_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2440__A1 (.DIODE(_0482_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2415__A1 (.DIODE(_0482_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2411__A1 (.DIODE(_0482_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2310__A1 (.DIODE(_0482_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2308__A1 (.DIODE(_0482_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2208__A (.DIODE(_0482_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3349__A1 (.DIODE(_0485_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2509__B (.DIODE(_0485_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2486__B (.DIODE(_0485_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2453__A (.DIODE(_0485_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2426__C1 (.DIODE(_0485_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2423__B (.DIODE(_0485_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2407__C (.DIODE(_0485_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2232__C1 (.DIODE(_0485_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2219__B (.DIODE(_0485_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2209__C1 (.DIODE(_0485_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3394__A1 (.DIODE(_0487_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3386__B2 (.DIODE(_0487_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3298__B1 (.DIODE(_0487_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2651__A2 (.DIODE(_0487_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2420__B (.DIODE(_0487_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2396__A1 (.DIODE(_0487_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2391__B (.DIODE(_0487_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2377__C (.DIODE(_0487_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2374__B (.DIODE(_0487_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2213__A (.DIODE(_0487_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3139__A1 (.DIODE(_0492_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3084__A0 (.DIODE(_0492_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3078__A1 (.DIODE(_0492_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2613__A (.DIODE(_0492_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2441__B (.DIODE(_0492_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2216__B (.DIODE(_0492_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2995__A1 (.DIODE(_0514_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2964__B (.DIODE(_0514_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2602__A (.DIODE(_0514_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2599__B1 (.DIODE(_0514_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2597__A1 (.DIODE(_0514_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2591__B1 (.DIODE(_0514_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2589__A (.DIODE(_0514_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2316__B (.DIODE(_0514_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2278__B2 (.DIODE(_0514_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2239__A (.DIODE(_0514_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3248__A2 (.DIODE(_0515_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3227__A2 (.DIODE(_0515_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3209__B2 (.DIODE(_0515_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3186__A2 (.DIODE(_0515_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3163__A2 (.DIODE(_0515_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3125__A2 (.DIODE(_0515_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2606__A2 (.DIODE(_0515_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2588__A2 (.DIODE(_0515_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2319__A2 (.DIODE(_0515_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2255__A2 (.DIODE(_0515_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4087__B (.DIODE(_0516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4083__B1 (.DIODE(_0516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2999__A (.DIODE(_0516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2988__B1 (.DIODE(_0516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2584__A (.DIODE(_0516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2363__B1 (.DIODE(_0516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2360__B (.DIODE(_0516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2253__B (.DIODE(_0516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3281__B2 (.DIODE(_0517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3125__A1 (.DIODE(_0517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3052__A0 (.DIODE(_0517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2751__B2 (.DIODE(_0517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2671__A1 (.DIODE(_0517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2669__A1 (.DIODE(_0517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2662__A (.DIODE(_0517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2321__A (.DIODE(_0517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2295__A (.DIODE(_0517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2252__B (.DIODE(_0517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3025__A3 (.DIODE(_0518_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3010__B (.DIODE(_0518_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2945__B (.DIODE(_0518_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2874__B (.DIODE(_0518_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2873__A (.DIODE(_0518_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2671__B1 (.DIODE(_0518_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2669__B1 (.DIODE(_0518_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2599__B2 (.DIODE(_0518_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2322__A (.DIODE(_0518_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2252__C (.DIODE(_0518_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3284__B2 (.DIODE(_0519_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3209__B1 (.DIODE(_0519_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2958__C (.DIODE(_0519_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2777__B2 (.DIODE(_0519_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2668__A1 (.DIODE(_0519_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2662__B (.DIODE(_0519_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2327__A (.DIODE(_0519_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2294__A (.DIODE(_0519_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2244__B (.DIODE(_0519_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3282__B2 (.DIODE(_0521_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3163__A1 (.DIODE(_0521_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3054__A0 (.DIODE(_0521_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2949__A1 (.DIODE(_0521_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2765__A2 (.DIODE(_0521_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2661__A (.DIODE(_0521_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2600__A (.DIODE(_0521_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2278__A1 (.DIODE(_0521_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2247__B2 (.DIODE(_0521_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2246__A1_N (.DIODE(_0521_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2289__A (.DIODE(_0530_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2255__B2 (.DIODE(_0530_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2668__A2 (.DIODE(_0551_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2662__C (.DIODE(_0551_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2277__B1 (.DIODE(_0551_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2964__C (.DIODE(_0576_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2858__C (.DIODE(_0576_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2667__B (.DIODE(_0576_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2313__A (.DIODE(_0576_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2858__D (.DIODE(_0585_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2667__C (.DIODE(_0585_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2312__D (.DIODE(_0585_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4086__A (.DIODE(_0589_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2989__A (.DIODE(_0589_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2965__A (.DIODE(_0589_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2795__A1 (.DIODE(_0589_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2747__A (.DIODE(_0589_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2654__A (.DIODE(_0589_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2595__A (.DIODE(_0589_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2578__A1 (.DIODE(_0589_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2362__A (.DIODE(_0589_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2316__A (.DIODE(_0589_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3280__B1 (.DIODE(_0591_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3002__A3 (.DIODE(_0591_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2997__B (.DIODE(_0591_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2606__B1 (.DIODE(_0591_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2599__A3 (.DIODE(_0591_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2598__A3 (.DIODE(_0591_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2590__A3 (.DIODE(_0591_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2588__B1 (.DIODE(_0591_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2365__A1 (.DIODE(_0591_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2318__C (.DIODE(_0591_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3072__B2 (.DIODE(_0597_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3021__A1 (.DIODE(_0597_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3010__A (.DIODE(_0597_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2960__A1 (.DIODE(_0597_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2946__A1 (.DIODE(_0597_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2874__A (.DIODE(_0597_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2859__A1 (.DIODE(_0597_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2593__A1 (.DIODE(_0597_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2585__A (.DIODE(_0597_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2354__A (.DIODE(_0597_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2586__C (.DIODE(_0626_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2354__C (.DIODE(_0626_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2959__C1 (.DIODE(_0631_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2787__B (.DIODE(_0631_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2779__C1 (.DIODE(_0631_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2359__C1 (.DIODE(_0631_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2636__A4 (.DIODE(_0634_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2364__A3 (.DIODE(_0634_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2363__A2 (.DIODE(_0634_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3331__A1 (.DIODE(_0641_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3220__A2 (.DIODE(_0641_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3205__A3 (.DIODE(_0641_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3202__B2 (.DIODE(_0641_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3132__B (.DIODE(_0641_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3131__A2 (.DIODE(_0641_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3129__A1 (.DIODE(_0641_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2370__D (.DIODE(_0641_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3064__B1 (.DIODE(_0644_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2649__A2 (.DIODE(_0644_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2392__B1 (.DIODE(_0644_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2388__A2 (.DIODE(_0644_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2379__A4 (.DIODE(_0644_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3408__A1 (.DIODE(_0652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3401__A1 (.DIODE(_0652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3395__S (.DIODE(_0652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3387__S (.DIODE(_0652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3072__A1 (.DIODE(_0652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2398__A1 (.DIODE(_0652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2396__B1 (.DIODE(_0652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2392__A1 (.DIODE(_0652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2383__A (.DIODE(_0652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2382__A (.DIODE(_0652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3351__A1 (.DIODE(_0678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2443__B (.DIODE(_0678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2411__A2 (.DIODE(_0678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3298__A2 (.DIODE(_0681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2610__A2 (.DIODE(_0681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2446__B (.DIODE(_0681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2432__B (.DIODE(_0681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2416__A (.DIODE(_0681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3122__A2 (.DIODE(_0709_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2451__B (.DIODE(_0709_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2444__C (.DIODE(_0709_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3220__A1 (.DIODE(_0760_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3197__B (.DIODE(_0760_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3170__A2 (.DIODE(_0760_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3168__A1 (.DIODE(_0760_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3166__A1 (.DIODE(_0760_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3142__A3 (.DIODE(_0760_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3140__A2 (.DIODE(_0760_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3131__A1 (.DIODE(_0760_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3088__C (.DIODE(_0760_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2496__B1 (.DIODE(_0760_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2826__B (.DIODE(_0780_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2823__A1 (.DIODE(_0780_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2819__B1 (.DIODE(_0780_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2814__A (.DIODE(_0780_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2805__A2 (.DIODE(_0780_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2799__A2 (.DIODE(_0780_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2774__A2 (.DIODE(_0780_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2768__A2 (.DIODE(_0780_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2759__A (.DIODE(_0780_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2526__A2 (.DIODE(_0780_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2913__S (.DIODE(_0826_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2911__S (.DIODE(_0826_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2905__A2 (.DIODE(_0826_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2847__B1 (.DIODE(_0826_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2845__A1_N (.DIODE(_0826_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2844__B (.DIODE(_0826_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2840__A3 (.DIODE(_0826_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2836__C (.DIODE(_0826_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2582__B2 (.DIODE(_0826_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2572__B1 (.DIODE(_0826_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3288__A2 (.DIODE(_0839_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3287__A2 (.DIODE(_0839_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3286__A2 (.DIODE(_0839_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3285__A2 (.DIODE(_0839_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3284__A2 (.DIODE(_0839_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3283__A2 (.DIODE(_0839_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3282__A2 (.DIODE(_0839_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3281__A2 (.DIODE(_0839_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3279__A2 (.DIODE(_0839_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2590__B1 (.DIODE(_0839_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3280__A2 (.DIODE(_0841_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3025__A4 (.DIODE(_0841_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2593__C1 (.DIODE(_0841_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3539__B (.DIODE(_0862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3305__A (.DIODE(_0862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2651__A3 (.DIODE(_0862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2624__A (.DIODE(_0862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2621__A (.DIODE(_0862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4179__B1 (.DIODE(_0951_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4167__A (.DIODE(_0951_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4081__B1 (.DIODE(_0951_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4078__C1 (.DIODE(_0951_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4071__B1 (.DIODE(_0951_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4065__B2 (.DIODE(_0951_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4040__A (.DIODE(_0951_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4037__A (.DIODE(_0951_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4009__A (.DIODE(_0951_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2744__A (.DIODE(_0951_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4085__A (.DIODE(_0979_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2959__A2 (.DIODE(_0979_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2808__A2 (.DIODE(_0979_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2779__A2 (.DIODE(_0979_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3020__A (.DIODE(_1054_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2994__A1 (.DIODE(_1054_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2869__B (.DIODE(_1054_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3565__B2 (.DIODE(_1119_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3523__A0 (.DIODE(_1119_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3486__A1 (.DIODE(_1119_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3443__A1 (.DIODE(_1119_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3424__A0 (.DIODE(_1119_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3352__B2 (.DIODE(_1119_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3309__A1 (.DIODE(_1119_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3290__A0 (.DIODE(_1119_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3281__A1 (.DIODE(_1119_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2967__A0 (.DIODE(_1119_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3054__S (.DIODE(_1122_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3052__S (.DIODE(_1122_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3050__S (.DIODE(_1122_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2985__S (.DIODE(_1122_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2982__S (.DIODE(_1122_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2979__S (.DIODE(_1122_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2976__S (.DIODE(_1122_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2973__S (.DIODE(_1122_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2970__S (.DIODE(_1122_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2967__S (.DIODE(_1122_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3566__B2 (.DIODE(_1124_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3525__A0 (.DIODE(_1124_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3488__A1 (.DIODE(_1124_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3445__A1 (.DIODE(_1124_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3426__A0 (.DIODE(_1124_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3353__B2 (.DIODE(_1124_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3311__A1 (.DIODE(_1124_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3292__A0 (.DIODE(_1124_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3282__A1 (.DIODE(_1124_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2970__A0 (.DIODE(_1124_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3578__A1 (.DIODE(_1126_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3567__B2 (.DIODE(_1126_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3527__A0 (.DIODE(_1126_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3490__A1 (.DIODE(_1126_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3447__A1 (.DIODE(_1126_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3428__A0 (.DIODE(_1126_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3354__B2 (.DIODE(_1126_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3313__A1 (.DIODE(_1126_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3283__A1 (.DIODE(_1126_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2973__A0 (.DIODE(_1126_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3580__A1 (.DIODE(_1128_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3568__B2 (.DIODE(_1128_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3529__A0 (.DIODE(_1128_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3492__A1 (.DIODE(_1128_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3449__A1 (.DIODE(_1128_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3430__A0 (.DIODE(_1128_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3355__B2 (.DIODE(_1128_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3315__A1 (.DIODE(_1128_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3284__A1 (.DIODE(_1128_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2976__A0 (.DIODE(_1128_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3582__A1 (.DIODE(_1130_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3569__B2 (.DIODE(_1130_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3531__A0 (.DIODE(_1130_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3494__A1 (.DIODE(_1130_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3451__A1 (.DIODE(_1130_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3432__A0 (.DIODE(_1130_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3356__B2 (.DIODE(_1130_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3317__A1 (.DIODE(_1130_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3285__A1 (.DIODE(_1130_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2979__A0 (.DIODE(_1130_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3570__B2 (.DIODE(_1132_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3533__A0 (.DIODE(_1132_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3496__A1 (.DIODE(_1132_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3453__A1 (.DIODE(_1132_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3434__A0 (.DIODE(_1132_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3361__A0 (.DIODE(_1132_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3357__B2 (.DIODE(_1132_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3319__A1 (.DIODE(_1132_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3286__A1 (.DIODE(_1132_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2982__A0 (.DIODE(_1132_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3571__B2 (.DIODE(_1134_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3535__A0 (.DIODE(_1134_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3516__A0 (.DIODE(_1134_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3481__A1 (.DIODE(_1134_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3455__A1 (.DIODE(_1134_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3436__A0 (.DIODE(_1134_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3358__B2 (.DIODE(_1134_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3321__A1 (.DIODE(_1134_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3287__A1 (.DIODE(_1134_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2985__A0 (.DIODE(_1134_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3572__B2 (.DIODE(_1171_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3537__A0 (.DIODE(_1171_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3518__A0 (.DIODE(_1171_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3483__A1 (.DIODE(_1171_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3457__A1 (.DIODE(_1171_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3438__A0 (.DIODE(_1171_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3359__A0 (.DIODE(_1171_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3296__A0 (.DIODE(_1171_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3288__A1 (.DIODE(_1171_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3050__A0 (.DIODE(_1171_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3266__A (.DIODE(_1220_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3258__A1 (.DIODE(_1220_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3256__A (.DIODE(_1220_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3254__A (.DIODE(_1220_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3155__A (.DIODE(_1220_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3119__B (.DIODE(_1220_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3118__A1 (.DIODE(_1220_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3117__A_N (.DIODE(_1220_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3113__A1 (.DIODE(_1220_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3106__A (.DIODE(_1220_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3658__B (.DIODE(_1221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3270__A (.DIODE(_1221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3238__A_N (.DIODE(_1221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3212__A_N (.DIODE(_1221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3192__A (.DIODE(_1221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3188__A (.DIODE(_1221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3176__A_N (.DIODE(_1221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3150__A_N (.DIODE(_1221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3146__A (.DIODE(_1221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3114__A1 (.DIODE(_1221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3257__S (.DIODE(_1222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3253__S (.DIODE(_1222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3241__S (.DIODE(_1222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3179__S (.DIODE(_1222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3156__S (.DIODE(_1222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3147__A (.DIODE(_1222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3119__A (.DIODE(_1222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3116__S (.DIODE(_1222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3110__S (.DIODE(_1222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3108__A (.DIODE(_1222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3269__S (.DIODE(_1223_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3265__S (.DIODE(_1223_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3237__S (.DIODE(_1223_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3215__S (.DIODE(_1223_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3211__S (.DIODE(_1223_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3187__S (.DIODE(_1223_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3175__S (.DIODE(_1223_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3149__S (.DIODE(_1223_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3115__S (.DIODE(_1223_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3109__S (.DIODE(_1223_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3663__C (.DIODE(_1227_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3272__B1 (.DIODE(_1227_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3243__B1 (.DIODE(_1227_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3217__B1 (.DIODE(_1227_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3194__B1 (.DIODE(_1227_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3181__B1 (.DIODE(_1227_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3158__B1 (.DIODE(_1227_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3151__A (.DIODE(_1227_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3118__C1 (.DIODE(_1227_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3113__B1 (.DIODE(_1227_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3122__B1 (.DIODE(_1236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3271__S (.DIODE(_1261_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3267__S (.DIODE(_1261_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3236__S (.DIODE(_1261_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3210__S (.DIODE(_1261_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3193__S (.DIODE(_1261_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3191__S (.DIODE(_1261_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3189__S (.DIODE(_1261_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3174__S (.DIODE(_1261_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3153__A (.DIODE(_1261_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3148__S (.DIODE(_1261_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3161__B1 (.DIODE(_1274_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3361__S (.DIODE(_1388_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3359__S (.DIODE(_1388_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3292__S (.DIODE(_1388_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3290__S (.DIODE(_1388_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3321__S (.DIODE(_1401_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3319__S (.DIODE(_1401_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3317__S (.DIODE(_1401_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3315__S (.DIODE(_1401_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3313__S (.DIODE(_1401_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3311__S (.DIODE(_1401_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3309__S (.DIODE(_1401_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3377__S (.DIODE(_1434_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3375__S (.DIODE(_1434_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3373__S (.DIODE(_1434_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3371__S (.DIODE(_1434_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3369__S (.DIODE(_1434_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3367__S (.DIODE(_1434_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3365__S (.DIODE(_1434_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3557__B (.DIODE(_1475_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3554__B (.DIODE(_1475_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3478__B (.DIODE(_1475_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3475__B (.DIODE(_1475_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3472__B (.DIODE(_1475_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3469__B (.DIODE(_1475_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3466__B (.DIODE(_1475_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3459__B (.DIODE(_1475_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3422__B (.DIODE(_1475_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3438__S (.DIODE(_1478_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3436__S (.DIODE(_1478_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3434__S (.DIODE(_1478_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3432__S (.DIODE(_1478_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3430__S (.DIODE(_1478_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3428__S (.DIODE(_1478_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3426__S (.DIODE(_1478_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3424__S (.DIODE(_1478_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3457__S (.DIODE(_1489_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3455__S (.DIODE(_1489_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3453__S (.DIODE(_1489_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3451__S (.DIODE(_1489_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3449__S (.DIODE(_1489_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3447__S (.DIODE(_1489_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3445__S (.DIODE(_1489_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3443__S (.DIODE(_1489_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3483__S (.DIODE(_1502_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3481__S (.DIODE(_1502_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3479__S (.DIODE(_1502_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3476__S (.DIODE(_1502_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3473__S (.DIODE(_1502_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3470__S (.DIODE(_1502_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3467__S (.DIODE(_1502_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3464__S (.DIODE(_1502_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3500__S (.DIODE(_1516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3498__S (.DIODE(_1516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3496__S (.DIODE(_1516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3494__S (.DIODE(_1516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3492__S (.DIODE(_1516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3490__S (.DIODE(_1516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3488__S (.DIODE(_1516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3486__S (.DIODE(_1516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3518__S (.DIODE(_1526_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3516__S (.DIODE(_1526_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3514__S (.DIODE(_1526_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3512__S (.DIODE(_1526_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3510__S (.DIODE(_1526_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3508__S (.DIODE(_1526_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3506__S (.DIODE(_1526_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3504__S (.DIODE(_1526_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3537__S (.DIODE(_1537_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3535__S (.DIODE(_1537_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3533__S (.DIODE(_1537_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3531__S (.DIODE(_1537_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3529__S (.DIODE(_1537_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3527__S (.DIODE(_1537_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3525__S (.DIODE(_1537_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3523__S (.DIODE(_1537_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3558__S (.DIODE(_1548_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3555__S (.DIODE(_1548_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3552__S (.DIODE(_1548_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3550__S (.DIODE(_1548_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3548__S (.DIODE(_1548_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3546__S (.DIODE(_1548_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3544__S (.DIODE(_1548_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3542__S (.DIODE(_1548_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3572__A2 (.DIODE(_1560_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3571__A2 (.DIODE(_1560_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3570__A2 (.DIODE(_1560_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3569__A2 (.DIODE(_1560_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3568__A2 (.DIODE(_1560_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3567__A2 (.DIODE(_1560_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3566__A2 (.DIODE(_1560_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3565__A2 (.DIODE(_1560_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3572__B1 (.DIODE(_1563_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3571__B1 (.DIODE(_1563_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3570__B1 (.DIODE(_1563_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3569__B1 (.DIODE(_1563_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3568__B1 (.DIODE(_1563_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3567__B1 (.DIODE(_1563_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3566__B1 (.DIODE(_1563_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3565__B1 (.DIODE(_1563_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3588__S (.DIODE(_1564_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3586__S (.DIODE(_1564_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3584__S (.DIODE(_1564_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3582__S (.DIODE(_1564_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3580__S (.DIODE(_1564_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3578__S (.DIODE(_1564_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3576__S (.DIODE(_1564_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3574__S (.DIODE(_1564_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4004__B1 (.DIODE(_1589_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4003__B (.DIODE(_1589_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3875__A_N (.DIODE(_1589_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3873__A_N (.DIODE(_1589_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3871__A_N (.DIODE(_1589_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3869__A_N (.DIODE(_1589_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3867__A_N (.DIODE(_1589_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3865__A_N (.DIODE(_1589_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3863__A_N (.DIODE(_1589_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3609__B (.DIODE(_1589_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3820__S (.DIODE(_1594_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3806__S (.DIODE(_1594_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3793__S (.DIODE(_1594_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3781__S (.DIODE(_1594_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3768__S (.DIODE(_1594_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3755__S (.DIODE(_1594_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3742__S (.DIODE(_1594_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3707__S (.DIODE(_1594_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3705__A (.DIODE(_1594_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3615__A (.DIODE(_1594_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3823__B_N (.DIODE(_1595_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3785__A1 (.DIODE(_1595_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3784__B_N (.DIODE(_1595_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3746__A1 (.DIODE(_1595_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3745__B_N (.DIODE(_1595_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3647__A1 (.DIODE(_1595_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3639__A (.DIODE(_1595_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3638__A (.DIODE(_1595_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3624__A1 (.DIODE(_1595_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3616__A (.DIODE(_1595_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3824__B1_N (.DIODE(_1598_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3811__A_N (.DIODE(_1598_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3798__A_N (.DIODE(_1598_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3785__B1_N (.DIODE(_1598_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3772__A_N (.DIODE(_1598_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3759__A_N (.DIODE(_1598_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3713__A (.DIODE(_1598_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3712__A_N (.DIODE(_1598_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3625__A (.DIODE(_1598_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3619__B (.DIODE(_1598_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3827__A2 (.DIODE(_1602_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3815__A2 (.DIODE(_1602_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3802__A2 (.DIODE(_1602_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3788__A2 (.DIODE(_1602_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3776__A2 (.DIODE(_1602_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3763__A2 (.DIODE(_1602_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3749__A2 (.DIODE(_1602_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3720__A2 (.DIODE(_1602_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3645__B1 (.DIODE(_1602_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3623__B (.DIODE(_1602_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3826__B2 (.DIODE(_1604_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3821__A_N (.DIODE(_1604_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3809__A1 (.DIODE(_1604_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3796__A1 (.DIODE(_1604_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3787__B2 (.DIODE(_1604_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3782__A_N (.DIODE(_1604_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3748__B2 (.DIODE(_1604_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3743__A_N (.DIODE(_1604_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3708__A_N (.DIODE(_1604_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3626__A (.DIODE(_1604_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3822__A1 (.DIODE(_1605_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3783__A1 (.DIODE(_1605_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3770__A1 (.DIODE(_1605_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3757__A1 (.DIODE(_1605_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3744__A1 (.DIODE(_1605_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3709__A1 (.DIODE(_1605_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3639__B (.DIODE(_1605_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3635__A1 (.DIODE(_1605_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3628__A (.DIODE(_1605_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3627__A (.DIODE(_1605_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3822__C1 (.DIODE(_1609_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3783__C1 (.DIODE(_1609_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3770__C1 (.DIODE(_1609_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3757__C1 (.DIODE(_1609_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3744__C1 (.DIODE(_1609_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3709__C1 (.DIODE(_1609_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3645__A1 (.DIODE(_1609_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3642__A1 (.DIODE(_1609_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3635__A2 (.DIODE(_1609_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3632__A (.DIODE(_1609_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3826__C1 (.DIODE(_1610_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3814__A1 (.DIODE(_1610_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3801__A1 (.DIODE(_1610_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3787__C1 (.DIODE(_1610_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3775__A1 (.DIODE(_1610_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3762__A1 (.DIODE(_1610_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3748__C1 (.DIODE(_1610_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3716__A1 (.DIODE(_1610_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3637__C (.DIODE(_1610_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3636__A1 (.DIODE(_1610_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3828__A1 (.DIODE(_1611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3814__B1 (.DIODE(_1611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3801__B1 (.DIODE(_1611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3789__A1 (.DIODE(_1611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3775__B1 (.DIODE(_1611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3762__B1 (.DIODE(_1611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3750__A1 (.DIODE(_1611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3716__B1 (.DIODE(_1611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3637__B (.DIODE(_1611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3636__A2 (.DIODE(_1611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3697__C (.DIODE(_1661_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3695__A2 (.DIODE(_1661_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4002__A2 (.DIODE(_1666_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4001__A1 (.DIODE(_1666_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4000__A1 (.DIODE(_1666_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3999__A1 (.DIODE(_1666_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3998__A1 (.DIODE(_1666_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3997__A1 (.DIODE(_1666_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3996__A1 (.DIODE(_1666_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3995__A1 (.DIODE(_1666_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3994__A1 (.DIODE(_1666_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3701__B1_N (.DIODE(_1666_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3825__S (.DIODE(_1670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3824__A1 (.DIODE(_1670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3819__S (.DIODE(_1670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3786__S (.DIODE(_1670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3780__S (.DIODE(_1670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3767__S (.DIODE(_1670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3754__S (.DIODE(_1670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3747__S (.DIODE(_1670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3741__S (.DIODE(_1670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3706__S (.DIODE(_1670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3812__S (.DIODE(_1675_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3807__S (.DIODE(_1675_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3799__S (.DIODE(_1675_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3794__S (.DIODE(_1675_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3773__S (.DIODE(_1675_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3771__S (.DIODE(_1675_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3760__S (.DIODE(_1675_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3758__S (.DIODE(_1675_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3714__S (.DIODE(_1675_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3711__S (.DIODE(_1675_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4077__B1 (.DIODE(_1684_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3827__B1 (.DIODE(_1684_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3815__C1 (.DIODE(_1684_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3802__C1 (.DIODE(_1684_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3788__B1 (.DIODE(_1684_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3776__C1 (.DIODE(_1684_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3763__C1 (.DIODE(_1684_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3749__B1 (.DIODE(_1684_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3730__B1 (.DIODE(_1684_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3720__C1 (.DIODE(_1684_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3902__B (.DIODE(_1790_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3899__B (.DIODE(_1790_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3896__B (.DIODE(_1790_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3893__B (.DIODE(_1790_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3890__B (.DIODE(_1790_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3887__B (.DIODE(_1790_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3884__B (.DIODE(_1790_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3879__B (.DIODE(_1790_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3854__A (.DIODE(_1790_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3835__A (.DIODE(_1790_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3851__S (.DIODE(_1792_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3849__S (.DIODE(_1792_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3847__S (.DIODE(_1792_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3845__S (.DIODE(_1792_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3843__S (.DIODE(_1792_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3841__S (.DIODE(_1792_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3839__S (.DIODE(_1792_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3837__S (.DIODE(_1792_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4001__A2 (.DIODE(_1806_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4000__A2 (.DIODE(_1806_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3999__A2 (.DIODE(_1806_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3998__A2 (.DIODE(_1806_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3997__A2 (.DIODE(_1806_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3996__A2 (.DIODE(_1806_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3995__A2 (.DIODE(_1806_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3994__A2 (.DIODE(_1806_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3924__B (.DIODE(_1806_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3861__A (.DIODE(_1806_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4004__A1 (.DIODE(_1810_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4002__A1 (.DIODE(_1810_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3990__A2 (.DIODE(_1810_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3989__A2 (.DIODE(_1810_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3988__A2 (.DIODE(_1810_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3987__A2 (.DIODE(_1810_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3986__A2 (.DIODE(_1810_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3985__A2 (.DIODE(_1810_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3984__A2 (.DIODE(_1810_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3863__B (.DIODE(_1810_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3903__S (.DIODE(_1821_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3900__S (.DIODE(_1821_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3897__S (.DIODE(_1821_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3894__S (.DIODE(_1821_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3891__S (.DIODE(_1821_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3888__S (.DIODE(_1821_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3885__S (.DIODE(_1821_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3882__S (.DIODE(_1821_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3922__S (.DIODE(_1839_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3920__S (.DIODE(_1839_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3918__S (.DIODE(_1839_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3916__S (.DIODE(_1839_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3914__S (.DIODE(_1839_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3912__S (.DIODE(_1839_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3910__S (.DIODE(_1839_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3908__S (.DIODE(_1839_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3940__S (.DIODE(_1849_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3938__S (.DIODE(_1849_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3936__S (.DIODE(_1849_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3934__S (.DIODE(_1849_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3932__S (.DIODE(_1849_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3930__S (.DIODE(_1849_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3928__S (.DIODE(_1849_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3926__S (.DIODE(_1849_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3959__S (.DIODE(_1860_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3957__S (.DIODE(_1860_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3955__S (.DIODE(_1860_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3953__S (.DIODE(_1860_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3951__S (.DIODE(_1860_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3949__S (.DIODE(_1860_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3947__S (.DIODE(_1860_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3945__S (.DIODE(_1860_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3978__S (.DIODE(_1871_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3976__S (.DIODE(_1871_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3974__S (.DIODE(_1871_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3972__S (.DIODE(_1871_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3970__S (.DIODE(_1871_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3968__S (.DIODE(_1871_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3966__S (.DIODE(_1871_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3964__S (.DIODE(_1871_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4175__C1 (.DIODE(_1891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4172__C1 (.DIODE(_1891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4154__C1 (.DIODE(_1891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4147__C1 (.DIODE(_1891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4106__C1 (.DIODE(_1891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4076__C1 (.DIODE(_1891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4073__A (.DIODE(_1891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4062__B (.DIODE(_1891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4022__A (.DIODE(_1891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4018__A (.DIODE(_1891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3071__B1 (.DIODE(_2003_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3022__A1 (.DIODE(_2003_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2996__A1 (.DIODE(_2003_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2876__A1 (.DIODE(_2003_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2803__A1 (.DIODE(_2003_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2636__B1 (.DIODE(_2003_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2591__A1 (.DIODE(_2003_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2360__A (.DIODE(_2003_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2252__A (.DIODE(_2003_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2093__A (.DIODE(_2003_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3393__A (.DIODE(_2006_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3384__A (.DIODE(_2006_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3323__A2 (.DIODE(_2006_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3100__A (.DIODE(_2006_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2992__B (.DIODE(_2006_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2510__A (.DIODE(_2006_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2385__A2 (.DIODE(_2006_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2220__B (.DIODE(_2006_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2219__A (.DIODE(_2006_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2167__A (.DIODE(_2006_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2864__A (.DIODE(_2007_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2619__B (.DIODE(_2007_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2356__B1 (.DIODE(_2007_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2137__B (.DIODE(_2007_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2096__B (.DIODE(_2007_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3325__A (.DIODE(_2009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3207__A1 (.DIODE(_2009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2664__A2 (.DIODE(_2009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2663__B (.DIODE(_2009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2419__A (.DIODE(_2009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2372__A (.DIODE(_2009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2211__A (.DIODE(_2009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2167__B (.DIODE(_2009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2143__B (.DIODE(_2009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2109__B (.DIODE(_2009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3327__B1 (.DIODE(_2020_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2484__A1 (.DIODE(_2020_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2419__B (.DIODE(_2020_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2380__B2 (.DIODE(_2020_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2197__B (.DIODE(_2020_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2109__C (.DIODE(_2020_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3249__B1_N (.DIODE(_2023_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3203__B (.DIODE(_2023_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3200__A1 (.DIODE(_2023_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3199__C1 (.DIODE(_2023_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3073__A (.DIODE(_2023_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2178__A (.DIODE(_2023_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2129__D (.DIODE(_2023_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2122__B (.DIODE(_2023_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2121__B (.DIODE(_2023_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2115__A_N (.DIODE(_2023_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2240__B (.DIODE(_2064_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2237__B (.DIODE(_2064_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2166__A3 (.DIODE(_2064_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3654__A2 (.DIODE(_2078_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3325__B (.DIODE(_2078_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2419__C (.DIODE(_2078_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2372__B (.DIODE(_2078_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2211__B (.DIODE(_2078_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2167__C (.DIODE(_2078_));
 sky130_fd_sc_hd__diode_2 ANTENNA_input1_A (.DIODE(io_in[17]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input2_A (.DIODE(io_in[18]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input3_A (.DIODE(io_in[19]));
 sky130_fd_sc_hd__diode_2 ANTENNA__4091__A (.DIODE(\usb2uart.u_uart.uart_rx_inst.m_axis_tdata_reg[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3984__A1 (.DIODE(\usb2uart.u_uart.uart_rx_inst.m_axis_tdata_reg[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3945__A1 (.DIODE(\usb2uart.u_uart.uart_rx_inst.m_axis_tdata_reg[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3908__A0 (.DIODE(\usb2uart.u_uart.uart_rx_inst.m_axis_tdata_reg[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3879__A (.DIODE(\usb2uart.u_uart.uart_rx_inst.m_axis_tdata_reg[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3863__C (.DIODE(\usb2uart.u_uart.uart_rx_inst.m_axis_tdata_reg[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3837__A0 (.DIODE(\usb2uart.u_uart.uart_rx_inst.m_axis_tdata_reg[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4093__A (.DIODE(\usb2uart.u_uart.uart_rx_inst.m_axis_tdata_reg[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3985__A1 (.DIODE(\usb2uart.u_uart.uart_rx_inst.m_axis_tdata_reg[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3947__A1 (.DIODE(\usb2uart.u_uart.uart_rx_inst.m_axis_tdata_reg[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3910__A0 (.DIODE(\usb2uart.u_uart.uart_rx_inst.m_axis_tdata_reg[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3884__A (.DIODE(\usb2uart.u_uart.uart_rx_inst.m_axis_tdata_reg[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3865__C (.DIODE(\usb2uart.u_uart.uart_rx_inst.m_axis_tdata_reg[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3839__A0 (.DIODE(\usb2uart.u_uart.uart_rx_inst.m_axis_tdata_reg[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4095__A (.DIODE(\usb2uart.u_uart.uart_rx_inst.m_axis_tdata_reg[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3986__A1 (.DIODE(\usb2uart.u_uart.uart_rx_inst.m_axis_tdata_reg[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3949__A1 (.DIODE(\usb2uart.u_uart.uart_rx_inst.m_axis_tdata_reg[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3912__A0 (.DIODE(\usb2uart.u_uart.uart_rx_inst.m_axis_tdata_reg[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3887__A (.DIODE(\usb2uart.u_uart.uart_rx_inst.m_axis_tdata_reg[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3867__C (.DIODE(\usb2uart.u_uart.uart_rx_inst.m_axis_tdata_reg[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3841__A0 (.DIODE(\usb2uart.u_uart.uart_rx_inst.m_axis_tdata_reg[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4099__A (.DIODE(\usb2uart.u_uart.uart_rx_inst.m_axis_tdata_reg[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3988__A1 (.DIODE(\usb2uart.u_uart.uart_rx_inst.m_axis_tdata_reg[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3953__A1 (.DIODE(\usb2uart.u_uart.uart_rx_inst.m_axis_tdata_reg[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3916__A0 (.DIODE(\usb2uart.u_uart.uart_rx_inst.m_axis_tdata_reg[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3893__A (.DIODE(\usb2uart.u_uart.uart_rx_inst.m_axis_tdata_reg[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3871__C (.DIODE(\usb2uart.u_uart.uart_rx_inst.m_axis_tdata_reg[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3845__A0 (.DIODE(\usb2uart.u_uart.uart_rx_inst.m_axis_tdata_reg[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4101__A (.DIODE(\usb2uart.u_uart.uart_rx_inst.m_axis_tdata_reg[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3989__A1 (.DIODE(\usb2uart.u_uart.uart_rx_inst.m_axis_tdata_reg[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3955__A1 (.DIODE(\usb2uart.u_uart.uart_rx_inst.m_axis_tdata_reg[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3918__A0 (.DIODE(\usb2uart.u_uart.uart_rx_inst.m_axis_tdata_reg[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3896__A (.DIODE(\usb2uart.u_uart.uart_rx_inst.m_axis_tdata_reg[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3873__C (.DIODE(\usb2uart.u_uart.uart_rx_inst.m_axis_tdata_reg[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3847__A0 (.DIODE(\usb2uart.u_uart.uart_rx_inst.m_axis_tdata_reg[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4103__A (.DIODE(\usb2uart.u_uart.uart_rx_inst.m_axis_tdata_reg[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3990__A1 (.DIODE(\usb2uart.u_uart.uart_rx_inst.m_axis_tdata_reg[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3957__A1 (.DIODE(\usb2uart.u_uart.uart_rx_inst.m_axis_tdata_reg[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3920__A0 (.DIODE(\usb2uart.u_uart.uart_rx_inst.m_axis_tdata_reg[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3899__A (.DIODE(\usb2uart.u_uart.uart_rx_inst.m_axis_tdata_reg[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3875__C (.DIODE(\usb2uart.u_uart.uart_rx_inst.m_axis_tdata_reg[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3849__A0 (.DIODE(\usb2uart.u_uart.uart_rx_inst.m_axis_tdata_reg[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4105__A (.DIODE(\usb2uart.u_uart.uart_rx_inst.m_axis_tdata_reg[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3991__A0 (.DIODE(\usb2uart.u_uart.uart_rx_inst.m_axis_tdata_reg[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3959__A1 (.DIODE(\usb2uart.u_uart.uart_rx_inst.m_axis_tdata_reg[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3922__A0 (.DIODE(\usb2uart.u_uart.uart_rx_inst.m_axis_tdata_reg[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3902__A (.DIODE(\usb2uart.u_uart.uart_rx_inst.m_axis_tdata_reg[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3878__A1 (.DIODE(\usb2uart.u_uart.uart_rx_inst.m_axis_tdata_reg[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3851__A0 (.DIODE(\usb2uart.u_uart.uart_rx_inst.m_axis_tdata_reg[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3405__S (.DIODE(\usb2uart.u_usb_cdc.bulk_out_nak ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3400__S (.DIODE(\usb2uart.u_usb_cdc.bulk_out_nak ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3391__S (.DIODE(\usb2uart.u_usb_cdc.bulk_out_nak ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3385__S (.DIODE(\usb2uart.u_usb_cdc.bulk_out_nak ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3306__B2 (.DIODE(\usb2uart.u_usb_cdc.bulk_out_nak ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2988__A2 (.DIODE(\usb2uart.u_usb_cdc.bulk_out_nak ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2956__A (.DIODE(\usb2uart.u_usb_cdc.bulk_out_nak ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3050__A1 (.DIODE(\usb2uart.u_usb_cdc.endp[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2871__A1 (.DIODE(\usb2uart.u_usb_cdc.endp[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2870__A1 (.DIODE(\usb2uart.u_usb_cdc.endp[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2862__S (.DIODE(\usb2uart.u_usb_cdc.endp[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2775__S (.DIODE(\usb2uart.u_usb_cdc.endp[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2652__A (.DIODE(\usb2uart.u_usb_cdc.endp[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2619__A (.DIODE(\usb2uart.u_usb_cdc.endp[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2137__A (.DIODE(\usb2uart.u_usb_cdc.endp[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2096__A_N (.DIODE(\usb2uart.u_usb_cdc.endp[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3674__A (.DIODE(\usb2uart.u_usb_cdc.in_data_ack ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2990__C_N (.DIODE(\usb2uart.u_usb_cdc.in_data_ack ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2876__B2 (.DIODE(\usb2uart.u_usb_cdc.in_data_ack ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2395__A2 (.DIODE(\usb2uart.u_usb_cdc.in_data_ack ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2394__A2 (.DIODE(\usb2uart.u_usb_cdc.in_data_ack ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2392__A2 (.DIODE(\usb2uart.u_usb_cdc.in_data_ack ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2376__A2 (.DIODE(\usb2uart.u_usb_cdc.in_data_ack ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2374__A (.DIODE(\usb2uart.u_usb_cdc.in_data_ack ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3469__A (.DIODE(\usb2uart.u_usb_cdc.out_data[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2972__A (.DIODE(\usb2uart.u_usb_cdc.out_data[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2452__A (.DIODE(\usb2uart.u_usb_cdc.out_data[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2447__A (.DIODE(\usb2uart.u_usb_cdc.out_data[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2310__B2 (.DIODE(\usb2uart.u_usb_cdc.out_data[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2305__A1 (.DIODE(\usb2uart.u_usb_cdc.out_data[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2284__A (.DIODE(\usb2uart.u_usb_cdc.out_data[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2282__A (.DIODE(\usb2uart.u_usb_cdc.out_data[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2206__A (.DIODE(\usb2uart.u_usb_cdc.out_data[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2193__A (.DIODE(\usb2uart.u_usb_cdc.out_data[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3472__A (.DIODE(\usb2uart.u_usb_cdc.out_data[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2975__A (.DIODE(\usb2uart.u_usb_cdc.out_data[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2305__B2 (.DIODE(\usb2uart.u_usb_cdc.out_data[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2288__B (.DIODE(\usb2uart.u_usb_cdc.out_data[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2206__B (.DIODE(\usb2uart.u_usb_cdc.out_data[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2192__A (.DIODE(\usb2uart.u_usb_cdc.out_data[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3475__A (.DIODE(\usb2uart.u_usb_cdc.out_data[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2978__A (.DIODE(\usb2uart.u_usb_cdc.out_data[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2444__A_N (.DIODE(\usb2uart.u_usb_cdc.out_data[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2440__B1 (.DIODE(\usb2uart.u_usb_cdc.out_data[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2414__A (.DIODE(\usb2uart.u_usb_cdc.out_data[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2307__A (.DIODE(\usb2uart.u_usb_cdc.out_data[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2290__A (.DIODE(\usb2uart.u_usb_cdc.out_data[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2281__B (.DIODE(\usb2uart.u_usb_cdc.out_data[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2190__A (.DIODE(\usb2uart.u_usb_cdc.out_data[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3584__A1 (.DIODE(\usb2uart.u_usb_cdc.out_data[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3478__A (.DIODE(\usb2uart.u_usb_cdc.out_data[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2981__A (.DIODE(\usb2uart.u_usb_cdc.out_data[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2443__D (.DIODE(\usb2uart.u_usb_cdc.out_data[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2309__A (.DIODE(\usb2uart.u_usb_cdc.out_data[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2284__B (.DIODE(\usb2uart.u_usb_cdc.out_data[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2190__B (.DIODE(\usb2uart.u_usb_cdc.out_data[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3588__A1 (.DIODE(\usb2uart.u_usb_cdc.out_data[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3557__A (.DIODE(\usb2uart.u_usb_cdc.out_data[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3500__A1 (.DIODE(\usb2uart.u_usb_cdc.out_data[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3307__A1 (.DIODE(\usb2uart.u_usb_cdc.out_data[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3049__A (.DIODE(\usb2uart.u_usb_cdc.out_data[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2478__A1 (.DIODE(\usb2uart.u_usb_cdc.out_data[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2410__A (.DIODE(\usb2uart.u_usb_cdc.out_data[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2282__B (.DIODE(\usb2uart.u_usb_cdc.out_data[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2214__A (.DIODE(\usb2uart.u_usb_cdc.out_data[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2191__A (.DIODE(\usb2uart.u_usb_cdc.out_data[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3810__S (.DIODE(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_first_q[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3797__S (.DIODE(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_first_q[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3710__A (.DIODE(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_first_q[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3619__A (.DIODE(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_first_q[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3614__A (.DIODE(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_first_q[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3592__B (.DIODE(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_first_q[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3809__C1 (.DIODE(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_first_q[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3796__C1 (.DIODE(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_first_q[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3631__A (.DIODE(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_first_q[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3620__A (.DIODE(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_first_q[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3594__B (.DIODE(\usb2uart.u_usb_cdc.u_bulk_endp.u_out_fifo.out_first_q[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3348__A1 (.DIODE(\usb2uart.u_usb_cdc.u_ctrl_endp.byte_cnt_q[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3347__A1 (.DIODE(\usb2uart.u_usb_cdc.u_ctrl_endp.byte_cnt_q[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3276__B1 (.DIODE(\usb2uart.u_usb_cdc.u_ctrl_endp.byte_cnt_q[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3205__B1 (.DIODE(\usb2uart.u_usb_cdc.u_ctrl_endp.byte_cnt_q[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3102__A_N (.DIODE(\usb2uart.u_usb_cdc.u_ctrl_endp.byte_cnt_q[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2178__C (.DIODE(\usb2uart.u_usb_cdc.u_ctrl_endp.byte_cnt_q[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2129__B_N (.DIODE(\usb2uart.u_usb_cdc.u_ctrl_endp.byte_cnt_q[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2125__B (.DIODE(\usb2uart.u_usb_cdc.u_ctrl_endp.byte_cnt_q[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2115__C (.DIODE(\usb2uart.u_usb_cdc.u_ctrl_endp.byte_cnt_q[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2104__C (.DIODE(\usb2uart.u_usb_cdc.u_ctrl_endp.byte_cnt_q[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3069__A0 (.DIODE(\usb2uart.u_usb_cdc.u_ctrl_endp.dev_state_qq[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2539__A2 (.DIODE(\usb2uart.u_usb_cdc.u_ctrl_endp.dev_state_qq[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2445__A2 (.DIODE(\usb2uart.u_usb_cdc.u_ctrl_endp.dev_state_qq[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2442__B (.DIODE(\usb2uart.u_usb_cdc.u_ctrl_endp.dev_state_qq[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2406__A2 (.DIODE(\usb2uart.u_usb_cdc.u_ctrl_endp.dev_state_qq[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2135__A2 (.DIODE(\usb2uart.u_usb_cdc.u_ctrl_endp.dev_state_qq[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2445__B1_N (.DIODE(\usb2uart.u_usb_cdc.u_ctrl_endp.in_dir_q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2406__B1 (.DIODE(\usb2uart.u_usb_cdc.u_ctrl_endp.in_dir_q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2184__A (.DIODE(\usb2uart.u_usb_cdc.u_ctrl_endp.in_dir_q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2102__D (.DIODE(\usb2uart.u_usb_cdc.u_ctrl_endp.in_dir_q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2098__A_N (.DIODE(\usb2uart.u_usb_cdc.u_ctrl_endp.in_dir_q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3122__A1 (.DIODE(\usb2uart.u_usb_cdc.u_ctrl_endp.req_q[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2630__B1 (.DIODE(\usb2uart.u_usb_cdc.u_ctrl_endp.req_q[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2476__A (.DIODE(\usb2uart.u_usb_cdc.u_ctrl_endp.req_q[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2471__A (.DIODE(\usb2uart.u_usb_cdc.u_ctrl_endp.req_q[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2436__A (.DIODE(\usb2uart.u_usb_cdc.u_ctrl_endp.req_q[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2228__A (.DIODE(\usb2uart.u_usb_cdc.u_ctrl_endp.req_q[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2132__A (.DIODE(\usb2uart.u_usb_cdc.u_ctrl_endp.req_q[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4083__A1 (.DIODE(\usb2uart.u_usb_cdc.u_ctrl_endp.req_q[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3298__A1 (.DIODE(\usb2uart.u_usb_cdc.u_ctrl_endp.req_q[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3068__A1 (.DIODE(\usb2uart.u_usb_cdc.u_ctrl_endp.req_q[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3061__A1 (.DIODE(\usb2uart.u_usb_cdc.u_ctrl_endp.req_q[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3059__A (.DIODE(\usb2uart.u_usb_cdc.u_ctrl_endp.req_q[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2993__A_N (.DIODE(\usb2uart.u_usb_cdc.u_ctrl_endp.req_q[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2504__B1 (.DIODE(\usb2uart.u_usb_cdc.u_ctrl_endp.req_q[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2477__A1 (.DIODE(\usb2uart.u_usb_cdc.u_ctrl_endp.req_q[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2469__A (.DIODE(\usb2uart.u_usb_cdc.u_ctrl_endp.req_q[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2435__B (.DIODE(\usb2uart.u_usb_cdc.u_ctrl_endp.req_q[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3283__B2 (.DIODE(\usb2uart.u_usb_cdc.u_sie.data_q[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3186__A1 (.DIODE(\usb2uart.u_usb_cdc.u_sie.data_q[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3056__A0 (.DIODE(\usb2uart.u_usb_cdc.u_sie.data_q[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2770__A2_N (.DIODE(\usb2uart.u_usb_cdc.u_sie.data_q[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2326__A (.DIODE(\usb2uart.u_usb_cdc.u_sie.data_q[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2286__A (.DIODE(\usb2uart.u_usb_cdc.u_sie.data_q[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2268__C1 (.DIODE(\usb2uart.u_usb_cdc.u_sie.data_q[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2250__A (.DIODE(\usb2uart.u_usb_cdc.u_sie.data_q[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2249__C_N (.DIODE(\usb2uart.u_usb_cdc.u_sie.data_q[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3285__B2 (.DIODE(\usb2uart.u_usb_cdc.u_sie.data_q[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3227__A1 (.DIODE(\usb2uart.u_usb_cdc.u_sie.data_q[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2785__B2 (.DIODE(\usb2uart.u_usb_cdc.u_sie.data_q[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2332__A (.DIODE(\usb2uart.u_usb_cdc.u_sie.data_q[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2292__A (.DIODE(\usb2uart.u_usb_cdc.u_sie.data_q[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2247__A2_N (.DIODE(\usb2uart.u_usb_cdc.u_sie.data_q[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2246__B1 (.DIODE(\usb2uart.u_usb_cdc.u_sie.data_q[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3286__B2 (.DIODE(\usb2uart.u_usb_cdc.u_sie.data_q[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3248__A1 (.DIODE(\usb2uart.u_usb_cdc.u_sie.data_q[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2793__A2_N (.DIODE(\usb2uart.u_usb_cdc.u_sie.data_q[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2331__A (.DIODE(\usb2uart.u_usb_cdc.u_sie.data_q[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2299__A (.DIODE(\usb2uart.u_usb_cdc.u_sie.data_q[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2247__B1 (.DIODE(\usb2uart.u_usb_cdc.u_sie.data_q[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2246__A2_N (.DIODE(\usb2uart.u_usb_cdc.u_sie.data_q[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3287__B2 (.DIODE(\usb2uart.u_usb_cdc.u_sie.data_q[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3263__A0 (.DIODE(\usb2uart.u_usb_cdc.u_sie.data_q[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2802__A2 (.DIODE(\usb2uart.u_usb_cdc.u_sie.data_q[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2329__A (.DIODE(\usb2uart.u_usb_cdc.u_sie.data_q[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2297__S (.DIODE(\usb2uart.u_usb_cdc.u_sie.data_q[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2250__C_N (.DIODE(\usb2uart.u_usb_cdc.u_sie.data_q[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2249__B (.DIODE(\usb2uart.u_usb_cdc.u_sie.data_q[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3288__B2 (.DIODE(\usb2uart.u_usb_cdc.u_sie.data_q[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3279__A1 (.DIODE(\usb2uart.u_usb_cdc.u_sie.data_q[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2806__A2_N (.DIODE(\usb2uart.u_usb_cdc.u_sie.data_q[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2325__A (.DIODE(\usb2uart.u_usb_cdc.u_sie.data_q[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2280__A (.DIODE(\usb2uart.u_usb_cdc.u_sie.data_q[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2244__A (.DIODE(\usb2uart.u_usb_cdc.u_sie.data_q[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2516__A (.DIODE(\usb2uart.u_usb_cdc.u_sie.rx_err ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2315__A (.DIODE(\usb2uart.u_usb_cdc.u_sie.rx_err ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2166__A1 (.DIODE(\usb2uart.u_usb_cdc.u_sie.rx_err ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2156__B1 (.DIODE(\usb2uart.u_usb_cdc.u_sie.rx_err ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2134__B (.DIODE(\usb2uart.u_usb_cdc.u_sie.rx_err ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2091__A (.DIODE(\usb2uart.u_usb_cdc.u_sie.rx_err ));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_user_clock2_A (.DIODE(user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA_input4_A (.DIODE(wb_rst_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4874__A (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__4268__D (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__4875__A (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__4260__D (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__4107__B (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA__4107__A (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__4068__B1 (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__4031__B1 (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__4026__A (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__4011__B1 (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__3737__A (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__2925__B1 (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__2743__A (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__2741__A (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA_output6_A (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__4873__A (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__2659__A (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__2539__C1 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__2537__B2 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__2527__A (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__2152__A (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__2088__A (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA_output10_A (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__4078__A1 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout19_A (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout20_A (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA__4354__RESET_B (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout21_A (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout15_A (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout18_A (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout30_A (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout31_A (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA__4185__RESET_B (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout25_A (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout27_A (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout26_A (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout41_A (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout42_A (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout39_A (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__4342__RESET_B (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__4249__SET_B (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__4196__SET_B (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__4242__RESET_B (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA__4320__RESET_B (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout50_A (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA__4340__RESET_B (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA__4308__RESET_B (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA__4307__RESET_B (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA__4324__RESET_B (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA__4326__RESET_B (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA__4346__RESET_B (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA__4332__RESET_B (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA__4321__RESET_B (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA__4318__RESET_B (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA__4317__RESET_B (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA__4325__RESET_B (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA__4319__RESET_B (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA__4246__SET_B (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA__4323__RESET_B (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout51_A (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout52_A (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout46_A (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout49_A (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__4533__RESET_B (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__4565__RESET_B (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout43_A (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout34_A (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout38_A (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout53_A (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout22_A (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout32_A (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA__4392__RESET_B (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout61_A (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__4337__RESET_B (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__4338__RESET_B (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout58_A (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__4228__CLK (.DIODE(clknet_leaf_4_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA__4226__CLK (.DIODE(clknet_leaf_4_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA__4224__CLK (.DIODE(clknet_leaf_4_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA__4363__CLK (.DIODE(clknet_leaf_4_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA__4386__CLK (.DIODE(clknet_leaf_4_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA__4353__CLK (.DIODE(clknet_leaf_4_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA__4359__CLK (.DIODE(clknet_leaf_4_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA__4350__CLK (.DIODE(clknet_leaf_4_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA__4354__CLK (.DIODE(clknet_leaf_4_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA__4351__CLK (.DIODE(clknet_leaf_4_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA__4352__CLK (.DIODE(clknet_leaf_4_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA__4355__CLK (.DIODE(clknet_leaf_4_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA__4338__CLK (.DIODE(clknet_leaf_4_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA__4360__CLK (.DIODE(clknet_leaf_4_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA__4337__CLK (.DIODE(clknet_leaf_4_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA__4358__CLK (.DIODE(clknet_leaf_4_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA__4230__CLK (.DIODE(clknet_leaf_4_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA__4229__CLK (.DIODE(clknet_leaf_4_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA__4201__CLK (.DIODE(clknet_leaf_15_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA__4204__CLK (.DIODE(clknet_leaf_15_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA__4274__CLK (.DIODE(clknet_leaf_15_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA__4279__CLK (.DIODE(clknet_leaf_15_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA__4278__CLK (.DIODE(clknet_leaf_15_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA__4188__CLK (.DIODE(clknet_leaf_15_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA__4298__CLK (.DIODE(clknet_leaf_15_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA__4297__CLK (.DIODE(clknet_leaf_15_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA__4295__CLK (.DIODE(clknet_leaf_15_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA__4272__CLK (.DIODE(clknet_leaf_15_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA__4296__CLK (.DIODE(clknet_leaf_15_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA__4275__CLK (.DIODE(clknet_leaf_15_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA__4277__CLK (.DIODE(clknet_leaf_15_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA__4276__CLK (.DIODE(clknet_leaf_15_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA__4273__CLK (.DIODE(clknet_leaf_15_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA__4244__CLK (.DIODE(clknet_leaf_15_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA__4330__CLK (.DIODE(clknet_leaf_15_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA__4327__CLK (.DIODE(clknet_leaf_15_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA__4534__CLK (.DIODE(clknet_leaf_31_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA__4532__CLK (.DIODE(clknet_leaf_31_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA__4526__CLK (.DIODE(clknet_leaf_31_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA__4522__CLK (.DIODE(clknet_leaf_31_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA__4524__CLK (.DIODE(clknet_leaf_31_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA__4523__CLK (.DIODE(clknet_leaf_31_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA__4555__CLK (.DIODE(clknet_leaf_31_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA__4572__CLK (.DIODE(clknet_leaf_31_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA__4539__CLK (.DIODE(clknet_leaf_31_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA__4558__CLK (.DIODE(clknet_leaf_31_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA__4554__CLK (.DIODE(clknet_leaf_31_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA__4542__CLK (.DIODE(clknet_leaf_31_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA__4540__CLK (.DIODE(clknet_leaf_31_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA__4548__CLK (.DIODE(clknet_leaf_31_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA__4547__CLK (.DIODE(clknet_leaf_31_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA__4545__CLK (.DIODE(clknet_leaf_31_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA__4401__CLK (.DIODE(clknet_leaf_32_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA__4394__CLK (.DIODE(clknet_leaf_32_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA__4395__CLK (.DIODE(clknet_leaf_32_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA__4397__CLK (.DIODE(clknet_leaf_32_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA__4370__CLK (.DIODE(clknet_leaf_32_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA__4361__CLK (.DIODE(clknet_leaf_32_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA__4369__CLK (.DIODE(clknet_leaf_32_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA__4371__CLK (.DIODE(clknet_leaf_32_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA__4372__CLK (.DIODE(clknet_leaf_32_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA__4396__CLK (.DIODE(clknet_leaf_32_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA__4531__CLK (.DIODE(clknet_leaf_32_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA__4493__CLK (.DIODE(clknet_leaf_32_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA__4206__CLK (.DIODE(clknet_leaf_32_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA__4400__CLK (.DIODE(clknet_leaf_32_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA__4492__CLK (.DIODE(clknet_leaf_32_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA__4399__CLK (.DIODE(clknet_leaf_32_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA__4466__CLK (.DIODE(clknet_leaf_37_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA__4471__CLK (.DIODE(clknet_leaf_37_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA__4455__CLK (.DIODE(clknet_leaf_37_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA__4438__CLK (.DIODE(clknet_leaf_37_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA__4463__CLK (.DIODE(clknet_leaf_37_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA__4439__CLK (.DIODE(clknet_leaf_37_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA__4497__CLK (.DIODE(clknet_leaf_37_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA__4470__CLK (.DIODE(clknet_leaf_37_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA__4468__CLK (.DIODE(clknet_leaf_37_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA__4498__CLK (.DIODE(clknet_leaf_37_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA__4469__CLK (.DIODE(clknet_leaf_37_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA__4445__CLK (.DIODE(clknet_leaf_37_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA__4446__CLK (.DIODE(clknet_leaf_37_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA__4460__CLK (.DIODE(clknet_leaf_37_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA__4444__CLK (.DIODE(clknet_leaf_37_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA__4437__CLK (.DIODE(clknet_leaf_37_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA__4436__CLK (.DIODE(clknet_leaf_37_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_3__f_user_clock2_A (.DIODE(clknet_0_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_2__f_user_clock2_A (.DIODE(clknet_0_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_1__f_user_clock2_A (.DIODE(clknet_0_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_0__f_user_clock2_A (.DIODE(clknet_0_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_37_user_clock2_A (.DIODE(clknet_2_0__leaf_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_36_user_clock2_A (.DIODE(clknet_2_0__leaf_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_35_user_clock2_A (.DIODE(clknet_2_0__leaf_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_34_user_clock2_A (.DIODE(clknet_2_0__leaf_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_33_user_clock2_A (.DIODE(clknet_2_0__leaf_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_5_user_clock2_A (.DIODE(clknet_2_0__leaf_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_3_user_clock2_A (.DIODE(clknet_2_0__leaf_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_2_user_clock2_A (.DIODE(clknet_2_0__leaf_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_1_user_clock2_A (.DIODE(clknet_2_0__leaf_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_0_user_clock2_A (.DIODE(clknet_2_0__leaf_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_13_user_clock2_A (.DIODE(clknet_2_1__leaf_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_12_user_clock2_A (.DIODE(clknet_2_1__leaf_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_11_user_clock2_A (.DIODE(clknet_2_1__leaf_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_10_user_clock2_A (.DIODE(clknet_2_1__leaf_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_9_user_clock2_A (.DIODE(clknet_2_1__leaf_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_8_user_clock2_A (.DIODE(clknet_2_1__leaf_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA__4348__CLK (.DIODE(clknet_2_1__leaf_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_6_user_clock2_A (.DIODE(clknet_2_1__leaf_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_4_user_clock2_A (.DIODE(clknet_2_1__leaf_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_32_user_clock2_A (.DIODE(clknet_2_2__leaf_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_31_user_clock2_A (.DIODE(clknet_2_2__leaf_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_30_user_clock2_A (.DIODE(clknet_2_2__leaf_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_29_user_clock2_A (.DIODE(clknet_2_2__leaf_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_28_user_clock2_A (.DIODE(clknet_2_2__leaf_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_27_user_clock2_A (.DIODE(clknet_2_2__leaf_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_26_user_clock2_A (.DIODE(clknet_2_2__leaf_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_25_user_clock2_A (.DIODE(clknet_2_2__leaf_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_opt_1_0_user_clock2_A (.DIODE(clknet_2_2__leaf_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_23_user_clock2_A (.DIODE(clknet_2_2__leaf_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_22_user_clock2_A (.DIODE(clknet_2_2__leaf_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_21_user_clock2_A (.DIODE(clknet_2_3__leaf_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_20_user_clock2_A (.DIODE(clknet_2_3__leaf_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_19_user_clock2_A (.DIODE(clknet_2_3__leaf_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_18_user_clock2_A (.DIODE(clknet_2_3__leaf_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_17_user_clock2_A (.DIODE(clknet_2_3__leaf_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_16_user_clock2_A (.DIODE(clknet_2_3__leaf_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_15_user_clock2_A (.DIODE(clknet_2_3__leaf_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_14_user_clock2_A (.DIODE(clknet_2_3__leaf_user_clock2));
 sky130_ef_sc_hd__decap_12 FILLER_0_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_262 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_397 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_428 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_455 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_464 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_482 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_510 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_565 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_596 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_623 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_632 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_650 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_678 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_682 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_686 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_726 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_767 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_771 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_782 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_794 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_817 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_830 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_838 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_848 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_857 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_866 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_875 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_884 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_902 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_911 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_930 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_934 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_938 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_958 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_965 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_986 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_997 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1014 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1021 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1028 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1042 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1049 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1056 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1070 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1077 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1084 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1098 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1105 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1112 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1126 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1133 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1140 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1154 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1161 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1168 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1182 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1186 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1190 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1210 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1217 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1226 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1238 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1249 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1266 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1273 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1280 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1289 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1294 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1301 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1308 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1317 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1322 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1329 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1336 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1345 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1350 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1357 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1364 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1373 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1378 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1385 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1392 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1401 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1406 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1413 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1420 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1429 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1434 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1438 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1442 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1451 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1455 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1457 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1462 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1469 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1478 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1485 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1490 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1501 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1511 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1513 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1518 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1525 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1532 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1541 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1546 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1553 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1560 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1569 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1574 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1581 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1588 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1597 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1602 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1609 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1616 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1625 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1630 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1637 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1644 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1653 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1658 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1665 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1672 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1681 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1686 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1690 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1694 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1703 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1707 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1714 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1726 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1749 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1777 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1805 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1833 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1861 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1889 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_536 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_704 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_716 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1157 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1172 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1401 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1424 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1436 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_1448 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1661 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1676 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1693 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1721 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_993 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_1029 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1055 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1067 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1079 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_965 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_977 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_995 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1018 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_1030 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_1041 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1045 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_1053 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_987 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_998 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1004 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_1013 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_1022 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_1028 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_1037 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_1047 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_1069 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_853 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_871 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_874 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_885 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_893 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_914 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_920 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_932 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_944 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_965 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_985 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_1001 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1031 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_1048 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_1058 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1069 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_1086 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1094 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1106 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_1118 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_837 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_851 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_874 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_973 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_978 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_1013 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_1021 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_1028 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_1046 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1053 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_1075 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_1083 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_1111 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1118 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1130 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_1142 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_839 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_865 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_873 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_883 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_906 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_912 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_920 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_930 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_969 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_986 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_994 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_1000 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_1006 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1015 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_1021 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_1030 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1038 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1042 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1091 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_1098 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1128 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1140 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1152 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1164 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_847 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_855 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_859 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_891 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_896 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_916 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_945 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_957 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_969 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_1012 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_1032 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_1055 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1075 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_1108 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1130 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_1142 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_839 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_863 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_883 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_895 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_908 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_926 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_938 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_953 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_972 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_992 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_1000 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_1015 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_1028 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1045 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_1074 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_1084 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_1091 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1099 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_1116 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_825 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_850 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_857 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_861 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_913 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_934 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_942 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_954 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_966 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_979 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_987 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_992 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1011 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_1018 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_1028 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_1042 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_1049 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_1069 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_1080 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_1090 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_1107 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1125 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_1137 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_825 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_828 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_859 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_868 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_874 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_880 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_884 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_902 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_906 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_923 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_930 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_971 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_983 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_990 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_994 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_999 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_1021 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1039 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_1046 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_1062 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_1084 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_1091 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_1104 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1139 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1151 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1163 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_698 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_714 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_726 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_738 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_761 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_773 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_784 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_790 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_810 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_825 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_845 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_874 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_880 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_884 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_933 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_941 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_960 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_968 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_978 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_994 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_1004 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_1015 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_1024 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_1048 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1055 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_1067 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_1079 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1085 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_1111 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1118 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1130 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_1142 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_653 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_670 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_681 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_695 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_698 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_706 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_747 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_753 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_759 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_767 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_773 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_779 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_782 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_801 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_804 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_828 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_847 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_856 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_865 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_871 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_906 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_919 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_922 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_928 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_934 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_944 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_969 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_974 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_986 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_995 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_1004 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_1019 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_1028 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_1048 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_1055 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_1061 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1089 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_1095 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_1105 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_1125 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1131 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_1143 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1153 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_1165 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_1173 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1181 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1193 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1217 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_641 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_662 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_668 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_674 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_680 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_686 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_713 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_717 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_735 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_774 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_780 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_786 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_792 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_832 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_836 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_840 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_848 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_858 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_865 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_876 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_885 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_894 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_902 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_952 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_960 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_972 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1007 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_1024 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_1032 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_1046 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_1052 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1060 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_1077 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_1088 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_1097 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_1120 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_1126 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_1132 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_1138 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_1144 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_1153 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_1163 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_1169 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_1175 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_1181 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_1187 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1191 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_1194 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_1200 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_1209 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_1216 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_1224 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1242 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_1254 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_639 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_648 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_654 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_670 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_682 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_702 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_749 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_759 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_772 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_816 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_823 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_827 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_859 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_870 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_883 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_911 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_918 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_940 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_950 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_972 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_980 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_984 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_991 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_1006 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1015 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_1032 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_1043 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_1074 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_1085 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_1097 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_1143 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_1155 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1161 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_1164 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_1182 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1190 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_1193 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_1199 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1213 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_1216 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_1222 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_1228 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_1237 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_1243 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_1249 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_1255 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1267 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_1279 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_616 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_628 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_642 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_660 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_724 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_746 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_754 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_776 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_798 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_811 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_839 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_846 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_890 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_898 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_904 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_916 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_921 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_925 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_939 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_951 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_956 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_962 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1003 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_1020 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_1055 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_1061 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_1083 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_1103 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_1109 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_1133 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_1142 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_1175 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1203 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_1205 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_1227 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_1242 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_1248 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1254 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_1258 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_1272 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1278 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1290 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1302 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_1314 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_630 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_670 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_756 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_790 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_798 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_808 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_816 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_839 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_847 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_865 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_874 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_902 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_906 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_929 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_938 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_960 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_967 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_971 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_1002 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_1065 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_1069 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1075 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_1084 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_1105 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_1111 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_1117 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_1126 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_1154 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_1163 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1175 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1181 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_1191 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1197 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_1201 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_1214 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_1220 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1226 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_1255 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_1279 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_596 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_608 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_632 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_656 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_672 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_733 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_764 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_774 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_827 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_844 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_857 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_866 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_892 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_901 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_908 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_914 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_935 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_943 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_951 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_955 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_972 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_988 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_994 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_1012 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_1024 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_1041 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1045 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_1062 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_1074 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_1080 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_1100 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_1107 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_1122 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_1135 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_1142 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_1160 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_1173 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_1179 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_1198 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_1217 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_1223 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_1229 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1237 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_1247 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1251 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_1258 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_1261 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1265 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_1275 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_1281 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_1287 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_1293 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1299 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_1311 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_642 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_666 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_696 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_700 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_703 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_751 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_766 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_772 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_796 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_830 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_859 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_885 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_904 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_912 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_959 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_984 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_990 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_994 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_997 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_1006 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_1015 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_1036 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1044 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_1062 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_1085 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_1091 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1097 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_1132 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_1138 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_1151 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_1157 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1163 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_1173 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_1200 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_1206 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_1230 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1237 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_1258 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_1286 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_1289 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_1293 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_1299 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_1305 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1311 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1323 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_1335 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_603 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_610 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_618 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_662 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_720 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_779 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_826 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_850 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_857 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_891 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_923 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_931 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_952 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_962 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_968 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_991 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_999 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_1016 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_1030 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_1044 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_1053 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_1066 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_1090 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1097 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_1157 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_1181 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_1192 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_1202 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_1214 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_1225 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_1231 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1237 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_1258 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_1270 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_1281 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1293 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_1303 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1315 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_1317 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_1321 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1327 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1339 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1351 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_1363 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_603 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_639 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_670 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_702 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_739 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_752 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_779 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_782 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_790 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_812 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_838 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_847 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_858 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_865 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_879 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_883 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_895 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_903 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_927 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_939 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_946 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_959 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_967 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_973 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_997 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_1015 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_1038 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_1065 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_1070 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1076 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_1086 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_1110 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_1116 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_1126 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1134 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_1144 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_1150 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1154 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_1161 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_1181 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_1192 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1196 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_1217 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1223 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_1242 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_1253 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_1259 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_1265 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_1271 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_1277 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_1286 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_1289 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_1311 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_1318 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_1324 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1330 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_1342 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_563 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_575 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_621 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_666 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_675 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_687 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_712 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_723 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_731 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_752 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_780 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_786 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_799 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_817 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_835 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_843 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_851 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_855 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_867 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_878 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_890 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_899 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_911 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_948 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_958 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_966 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_970 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_976 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_991 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_998 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1004 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_1014 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_1024 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_1030 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_1037 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_1041 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_1067 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_1080 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_1104 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_1130 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1147 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_1158 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_1169 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_1175 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_1181 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_1194 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_1200 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_1205 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_1214 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1222 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_1243 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_1249 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1253 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_1257 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_1261 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_1272 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_1300 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_1308 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_1314 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_1317 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_1328 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1334 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1346 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1358 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_1370 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_541 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_639 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_650 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_658 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_694 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_704 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_744 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_863 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_872 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_883 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_894 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_932 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_938 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_962 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_1013 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_1039 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_1052 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_1058 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_1065 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_1076 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_1102 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_1108 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1112 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_1116 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_1132 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_1138 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1142 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_1163 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_1170 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_1188 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_1212 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_1222 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_1229 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_1233 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_1244 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1250 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_1271 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_1282 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_1289 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_1304 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_1332 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_1338 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1349 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1361 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1385 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_600 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_652 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_676 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_688 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_706 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_830 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_878 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_888 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_892 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_898 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_905 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_911 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_934 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_938 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_941 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_952 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_966 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_996 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_1020 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1024 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_1028 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_1048 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_1055 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_1068 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_1077 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_1086 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_1098 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_1105 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_1111 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_1117 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_1130 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_1137 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1147 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_1162 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_1168 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_1178 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_1184 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_1190 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_1202 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_1209 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_1215 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1223 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_1229 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_1243 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1247 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_1257 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_1261 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1267 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_1272 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1276 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_1284 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1290 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_1297 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1301 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_1308 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_1314 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_1317 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_1328 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_1335 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_1341 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_1347 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_1353 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1359 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_646 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_650 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_726 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_734 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_747 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_771 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_855 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_879 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_901 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_907 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_913 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_934 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_940 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_946 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_991 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_997 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_1020 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1028 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_1049 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_1055 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_1087 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_1111 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_1121 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_1132 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1138 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_1143 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_1156 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1164 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_1173 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1181 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_1202 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_1208 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1216 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_1226 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_1233 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_1238 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1244 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_1265 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_1276 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_1284 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_1289 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_1311 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_1335 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_1342 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_1345 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_1349 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_1355 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1361 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1385 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_620 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_626 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_662 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_698 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_707 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_734 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_767 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_795 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_820 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_828 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_842 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_867 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_892 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_915 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_929 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_936 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_942 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_966 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_972 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_976 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_985 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_1013 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1019 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_1022 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_1028 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_1034 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1041 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_1051 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_1075 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_1084 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_1104 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1108 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_1113 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_1125 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_1133 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1137 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_1154 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_1180 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_1186 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1190 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1203 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1211 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_1232 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_1242 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_1251 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_1257 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_1261 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_1275 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_1301 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_1314 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_1317 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_1332 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_1338 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_1344 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_1350 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_1356 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_1362 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_1368 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_632 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_670 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_688 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_766 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_804 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_814 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_848 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_859 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_867 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_878 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_938 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_946 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_964 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_970 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_991 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_997 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_1019 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_1028 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_1050 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1058 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_1065 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_1076 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1082 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_1103 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_1130 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_1140 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_1147 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_1153 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_1159 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1175 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_1184 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_1192 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_1203 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_1214 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1231 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_1240 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_1249 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_1259 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_1283 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1287 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_1289 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_1311 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1321 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_1342 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_1345 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_1349 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_1355 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1361 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1385 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_562 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_602 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_632 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_660 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_666 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_690 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_712 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_736 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_768 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_772 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_776 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_800 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_824 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_834 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_840 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_846 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_855 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_874 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_890 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_896 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_900 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_904 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_923 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_938 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_955 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_965 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_992 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_1018 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_1027 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_1033 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_1050 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_1056 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_1069 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_1075 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_1081 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_1104 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_1110 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_1120 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_1130 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1134 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_1144 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1155 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_1176 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1182 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_1202 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1209 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_1214 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_1223 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1229 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_1238 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_1252 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_1258 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_1261 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1265 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_1275 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_1286 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_1301 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_1314 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_1317 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_1321 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1325 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_1329 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_1335 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_1341 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_1347 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_1353 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_1359 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_534 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_583 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_628 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_680 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_708 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_736 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_770 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_796 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_824 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_838 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_850 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_863 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_870 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_922 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_935 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_941 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_964 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_974 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_983 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_999 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_1019 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_1025 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1029 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_1050 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1063 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1069 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_1090 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_1102 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1106 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_1121 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_1127 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_1153 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_1159 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1165 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_1172 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1181 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_1190 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1196 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_1217 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_1229 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_1255 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_1274 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1278 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_1286 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_1289 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1293 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_1303 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_1329 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_1335 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_1341 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_1345 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_1349 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_1355 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1361 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1385 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_513 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_562 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_630 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_656 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_663 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_675 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_688 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_730 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_773 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_794 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_800 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_834 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_838 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_846 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_876 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_888 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_945 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_952 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_962 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_1003 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1017 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_1027 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_1033 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_1049 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1053 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_1074 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_1082 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_1088 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_1103 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_1112 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_1123 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_1133 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1141 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_1160 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_1172 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1178 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1203 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_1205 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_1216 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_1231 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_1244 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1259 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_1261 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_1283 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1315 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_1317 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_1343 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_1349 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1355 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_1367 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_534 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_648 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_682 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_706 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_724 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_748 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_752 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_758 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_766 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_802 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_805 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_824 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_828 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_861 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_868 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_872 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_882 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_903 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_916 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_926 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_935 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_939 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_949 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_970 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_994 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_1031 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_1044 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_1052 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1058 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_1076 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1084 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_1105 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_1117 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_1125 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_1132 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_1145 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_1173 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_1199 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_1206 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_1216 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_1228 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_1241 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_1248 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_1259 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_1269 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_1278 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_1285 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_1289 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_1304 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_1311 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1319 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_1329 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_1336 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_1342 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_1345 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_1350 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1356 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1368 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1380 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_1392 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_513 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_616 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_626 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_661 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_672 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_705 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_715 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_736 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_762 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_770 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_824 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_828 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_831 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_850 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_867 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_873 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_922 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_934 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_944 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_950 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_959 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_968 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_978 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_987 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_1011 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_1023 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1029 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_1048 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1052 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_1062 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1066 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_1073 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_1079 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_1103 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1111 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_1132 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_1145 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_1155 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_1183 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_1195 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_1201 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_1205 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_1209 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_1221 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_1231 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1251 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_1258 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_1265 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_1289 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_1299 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_1314 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_1317 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1349 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_1361 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_568 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_592 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_623 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_630 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_670 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_686 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_690 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_694 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_702 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_708 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_714 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_740 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_744 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_792 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_816 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_838 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_847 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_864 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_871 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_880 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_907 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_911 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_919 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_922 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_930 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_939 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_949 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_974 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_1032 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_1056 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_1076 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_1100 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_1112 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_1132 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_1143 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_1159 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1165 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_1181 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_1187 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_1196 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_1209 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1213 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_1217 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_1239 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_1260 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1264 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_1273 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_1286 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_1289 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_1300 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1308 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_1318 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_1331 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_1341 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_1345 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_1349 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1355 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1367 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1379 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_1391 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_554 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_560 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_578 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_604 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_620 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_641 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_674 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_684 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_697 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_706 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_722 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_765 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_835 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_878 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_902 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_922 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_932 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_943 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_951 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_955 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_958 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_967 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_1004 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1035 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_1063 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_1072 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_1078 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_1084 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_1115 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_1122 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_1134 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_1144 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_1160 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_1169 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1181 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_1202 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_1214 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_1226 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1232 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_1241 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_1251 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_1258 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_1269 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1273 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_1277 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_1301 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_1314 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_1317 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_1321 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1351 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_1363 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_638 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_659 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_726 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_734 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_740 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_753 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_768 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_776 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_802 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_805 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_812 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_838 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_845 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_853 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_879 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_919 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_930 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_936 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_984 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_990 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_996 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1000 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1007 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1015 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_1029 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_1036 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1040 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_1044 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1048 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_1052 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_1069 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_1075 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_1099 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_1111 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_1131 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1135 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_1156 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_1166 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1170 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_1184 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_1190 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1196 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_1219 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_1229 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_1238 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_1265 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_1278 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_1286 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_1289 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_1297 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1301 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_1322 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_1329 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_1336 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_562 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_600 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_618 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_650 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_676 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_698 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_762 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_766 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_770 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_794 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_842 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_878 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_891 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_913 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_933 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_939 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_960 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_969 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_973 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_976 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_996 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_1002 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_1011 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_1027 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_1059 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_1065 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_1077 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_1086 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1099 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_1108 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_1132 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1136 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_1154 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_1160 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_1166 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_1182 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_1188 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1192 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_1201 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_1209 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_1236 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1242 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_1248 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_1257 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_1261 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1265 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_1286 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_1294 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_1302 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1315 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_1317 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_1328 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1334 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1346 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1358 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_1370 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_644 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_650 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_734 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_740 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_822 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_826 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_829 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_845 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_870 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_894 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_904 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_915 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_927 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_936 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_963 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_971 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_977 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_987 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_1000 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_1014 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_1024 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_1035 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_1046 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_1090 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_1096 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_1102 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_1108 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_1114 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_1125 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_1131 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_1144 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_1150 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_1177 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_1182 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1188 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_1196 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_1207 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1211 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_1218 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_1239 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_1266 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_1274 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1287 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_1289 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_1311 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_1318 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_1324 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1330 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_1342 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_562 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_618 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_684 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_768 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_772 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_781 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_824 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_830 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_890 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_896 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_902 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_908 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_932 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_942 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_948 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_959 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_978 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_988 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_1002 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_1013 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1019 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_1028 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_1037 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_1046 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_1055 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_1061 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_1067 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1071 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_1078 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_1099 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_1128 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1134 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_1142 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_1153 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1159 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_1163 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_1174 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_1180 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_1186 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1190 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_1198 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_1213 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_1219 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_1225 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_1231 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1235 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_1241 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_1248 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_1254 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_1265 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_1289 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_1295 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_1301 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_1307 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_559 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_590 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_596 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_628 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_670 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_678 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_702 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_746 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_782 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_790 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_800 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_835 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_850 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_858 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_882 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_888 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_919 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_936 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_960 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_967 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_983 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_994 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_1014 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1020 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_1024 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_1034 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_1044 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_1052 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_1062 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_1075 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_1083 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1087 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_1109 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1119 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1125 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_1140 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_1155 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_1170 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_1177 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_1188 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1194 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_1202 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_1209 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_1215 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1219 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1231 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_1243 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_1270 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1278 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_1282 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1293 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1305 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1329 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_557 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_586 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_618 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_650 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_667 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_672 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_680 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_707 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_715 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_724 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_730 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_776 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_780 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_783 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_794 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_810 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_827 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_830 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_837 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_848 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_866 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_904 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_908 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_912 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_947 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_959 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_969 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_999 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_1007 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_1014 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1027 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_1042 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_1054 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_1062 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_1077 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_1099 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1109 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_1130 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1138 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_1159 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1165 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_1175 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_1188 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1203 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_1216 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_1222 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_1228 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_1234 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_1240 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_1246 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_1252 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_1258 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_1269 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_1275 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1281 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1293 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_1305 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_590 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_596 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_614 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_631 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_644 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_702 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_736 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_742 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_749 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_761 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_768 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_794 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_800 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_808 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_814 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_845 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_858 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_864 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_872 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_883 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_907 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_911 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_917 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_926 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_932 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_940 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_957 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_969 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_975 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_990 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_1002 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_1019 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_1026 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1030 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_1038 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_1048 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_1062 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_1073 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_1081 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_1087 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_1097 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_1105 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_1132 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_1138 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_1144 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_1157 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_1163 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1167 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1175 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_1177 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_1181 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1187 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_1191 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1195 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_1201 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1207 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_1215 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_1223 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_1242 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_1248 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1254 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_1259 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_1266 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1272 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_1284 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_557 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_675 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_706 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_720 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_728 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_735 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_743 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_764 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_780 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_791 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_822 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_833 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_866 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_902 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_930 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_938 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_962 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_969 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_985 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_997 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_1004 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1010 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_1015 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1023 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_1032 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_1042 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_1048 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1056 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_1061 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_1072 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_1078 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_1103 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_1109 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1115 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_1119 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1125 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_1135 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_1142 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_1171 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_1184 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1192 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_1198 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_1205 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_1214 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_1223 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_1234 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_1244 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_1250 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_1258 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_590 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_596 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_614 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_632 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_636 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_679 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_683 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_805 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_814 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_848 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_855 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_866 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_877 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_888 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_894 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_905 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_913 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_917 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_924 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_943 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_962 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_972 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_979 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_990 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_1018 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_1028 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_1035 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_1041 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_1045 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_1075 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_1081 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_1087 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_1096 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_1102 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_1108 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_1114 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_1144 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_1151 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_1158 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_1164 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_1170 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_1199 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_1210 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_1220 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_1226 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_1243 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1273 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_557 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_667 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_675 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_708 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_723 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_735 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_775 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_786 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_792 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_824 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_828 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_834 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_846 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_857 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_890 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_906 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_913 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_938 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_947 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_966 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_985 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_1001 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_1024 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_1034 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_1045 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_1055 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_1063 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_1067 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_1075 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_1081 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_1125 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_1131 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_1157 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_1183 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_1189 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_1195 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_1201 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_1209 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1215 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1227 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1239 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_1251 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_580 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_637 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_643 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_662 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_700 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_706 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_749 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_759 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_792 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_799 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_810 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_839 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_850 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_859 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_868 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_876 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_887 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_894 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_912 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_920 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_941 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_958 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_962 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_966 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_970 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_979 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_991 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_1002 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_1014 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_1026 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_1038 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_1049 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_1058 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_1073 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1077 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_1084 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_1096 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_1102 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_1108 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1112 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_1116 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_1128 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_1134 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_1159 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1165 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_1181 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_1187 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_1193 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1199 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1211 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_1223 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_562 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_586 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_674 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_706 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_718 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_734 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_766 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_774 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_782 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_791 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_797 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_826 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_835 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_846 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_858 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_874 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_885 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_891 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_911 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_921 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_938 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_944 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_955 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_971 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_986 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_1005 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_1012 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_1023 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_1047 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_1055 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_1067 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_1083 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_1097 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1105 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_1113 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_1123 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_1132 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_1153 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_1159 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_1165 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_1171 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_1183 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_1189 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_1195 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_581 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_588 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_646 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_670 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_708 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_718 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_734 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_743 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_767 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_782 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_807 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_820 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_850 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_856 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_864 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_881 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_904 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_917 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_926 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_938 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_960 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_964 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_971 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_983 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_996 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_1016 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_1022 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_1034 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_1046 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_1062 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1071 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_1080 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_1092 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_1103 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1107 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_1111 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_1127 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_1133 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1137 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_1141 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_1147 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_1153 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_1159 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_1165 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1175 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_1181 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1187 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1199 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1211 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_1223 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_650 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_672 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_718 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_724 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_732 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_742 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_762 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_773 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_779 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_788 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_825 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_834 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_867 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_882 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_886 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_892 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_912 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_933 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_937 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_944 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_950 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_967 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_987 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_999 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_1012 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_1024 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_1028 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_1051 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_1065 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_1073 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_1079 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_1088 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_1117 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_1123 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_1144 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_1153 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_1159 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_1180 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1186 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_1198 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_541 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_578 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_602 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_670 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_791 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_820 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_838 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_850 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_861 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_870 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_879 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_887 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_894 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_915 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_951 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_964 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_970 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_982 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_990 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_997 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1007 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_1021 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_1047 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_1062 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1069 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_1075 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1079 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_1103 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1109 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_1117 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_1129 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_1137 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_1143 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_1155 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_1161 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_1167 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_1173 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1181 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1193 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1217 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_586 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_612 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_656 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_680 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_706 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_717 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_741 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_777 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_784 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_788 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_792 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_826 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_839 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_842 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_855 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_866 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_891 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_899 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_923 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_935 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_962 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_978 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_987 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_1008 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_1014 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_1023 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_1029 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_1033 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_1044 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_1050 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_1080 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_1098 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_1124 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_1136 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_1153 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_1183 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1189 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_610 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_623 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_639 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_648 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_705 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_762 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_794 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_800 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_803 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_815 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_852 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_860 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_870 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_894 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_922 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_933 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_940 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_958 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_969 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_1006 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1013 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_1034 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_1040 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1044 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_1065 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_1070 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_1083 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1097 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_1102 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_1109 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_1116 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_1135 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_1143 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_1150 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1156 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_1163 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1175 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_1181 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_1187 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_1193 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1199 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1211 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_1223 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_557 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_574 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_630 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_666 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_688 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_698 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_710 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_763 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_784 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_790 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_824 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_832 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_877 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_905 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_912 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_922 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_969 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_976 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_995 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_1005 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_1011 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_1015 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_1024 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_1062 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_1069 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_1075 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_1115 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_1125 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_1130 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_1137 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_1144 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_1171 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_1183 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_1189 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_1195 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_1201 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1209 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1221 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1245 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_646 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_683 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_687 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_696 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_702 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_708 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_778 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_812 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_837 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_847 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_868 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_876 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_884 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_895 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_958 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_964 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_968 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_972 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_976 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_984 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_996 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_1016 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_1022 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_1028 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_1041 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_1052 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_1076 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_1091 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_1116 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_1146 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_1173 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_1181 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_1187 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_1193 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_1199 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1211 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_1223 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_607 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_654 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_660 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_674 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_680 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_686 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_697 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_738 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_742 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_779 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_794 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_807 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_818 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_888 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_900 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_913 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_934 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_942 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_950 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_971 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_992 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_1004 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_1010 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_1020 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_1027 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_1037 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_1045 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_1051 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_1058 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_1071 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_1077 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_1097 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_1124 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_1130 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_1136 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_1142 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_1154 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_1160 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_1166 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_1172 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_1178 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_1202 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_1209 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_1215 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1221 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_1237 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1245 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_591 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_623 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_650 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_695 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_706 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_726 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_743 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_773 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_779 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_789 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_824 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_858 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_864 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_874 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_882 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_888 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_894 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_931 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_940 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_963 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_974 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_997 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1001 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_1006 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_1016 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_1027 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_1054 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_1060 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_1069 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1073 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_1081 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_1106 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_1112 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_1130 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_1140 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_1164 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_1170 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_1177 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_1181 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1187 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_1195 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_1201 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1231 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_1233 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_1242 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_1250 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1274 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_1286 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_616 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_656 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_676 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_695 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_716 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_726 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_753 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_763 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_777 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_801 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_824 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_828 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_856 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_866 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_879 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_888 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_896 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_902 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_910 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_934 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_941 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_945 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_964 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_968 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_971 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_990 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_997 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_1003 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_1013 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1027 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_1045 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1055 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_1076 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_1101 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_1126 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_1142 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_1164 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_1181 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_1192 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_1198 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_1214 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_1224 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_1230 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1234 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1242 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1254 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_1258 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1270 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1282 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1294 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_1306 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_1314 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_581 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_647 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_660 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_684 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_703 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_738 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_742 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_758 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_764 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_770 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_794 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_800 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_810 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_814 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_863 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_876 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_887 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_905 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_911 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_914 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_922 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_942 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_946 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_962 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_969 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_973 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_979 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_995 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_1031 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_1048 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_1052 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_1060 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_1073 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_1079 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_1091 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_1103 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_1129 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_1141 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_1158 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_1165 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_1175 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_1183 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_1197 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_1208 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_1218 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_1228 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_1237 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_1243 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_1247 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_1251 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_1259 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_1267 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1273 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_587 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_604 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_664 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_708 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_719 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_732 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_764 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_799 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_806 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_834 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_846 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_856 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_877 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_887 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_899 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_910 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_933 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_947 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_957 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_966 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_990 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_997 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1001 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1013 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_1020 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1028 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_1034 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1041 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_1049 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1053 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_1082 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_1088 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_1102 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_1110 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_1116 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1120 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_1129 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_1144 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1155 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_1176 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_1182 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_1193 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1203 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_1218 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_1229 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_1244 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_1251 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_1257 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1299 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_1311 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_585 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_634 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_682 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_686 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_708 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_723 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_738 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_749 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_766 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_778 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_812 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_836 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_847 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_868 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_879 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_883 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_916 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_936 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_940 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_946 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_969 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_976 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_980 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_995 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_999 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_1019 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_1025 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_1038 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1044 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_1051 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_1071 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_1082 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_1099 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1113 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_1117 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1127 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1143 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_1152 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_1158 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_1184 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_1191 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_1211 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_1221 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1231 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_1242 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1250 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_1258 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_1282 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_605 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_608 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_650 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_662 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_668 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_674 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_680 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_686 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_698 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_711 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_722 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_735 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_742 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_776 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_786 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_794 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_807 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_817 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_855 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_888 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_898 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_902 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_922 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_938 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_947 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_958 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_964 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_968 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_996 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_1017 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_1045 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_1053 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_1071 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_1081 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_1107 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_1113 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_1127 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_1138 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_1145 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_1159 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_1176 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_1183 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_1200 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_1209 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_1220 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_1226 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_1232 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_1258 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_1268 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1275 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1299 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_1311 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_625 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_631 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_652 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_658 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_696 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_702 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_708 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_726 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_749 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_760 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_779 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_818 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_847 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_856 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_864 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_885 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_935 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_946 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_977 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_992 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_996 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_1018 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_1024 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_1034 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_1055 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_1073 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_1079 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_1092 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_1099 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_1103 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_1112 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_1131 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_1147 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_1161 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_1168 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_1192 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_1200 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_1219 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_1231 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_1242 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_1253 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1270 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_1282 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_632 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_668 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_672 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_676 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_698 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_706 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_724 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_730 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_736 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_742 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_754 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_762 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_774 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_831 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_837 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_843 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_863 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_866 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_900 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_912 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_957 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_978 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_995 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_1022 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1028 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_1044 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_1068 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_1075 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1079 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_1100 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_1113 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_1124 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_1135 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_1158 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_1164 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_1188 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1194 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_1202 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_1205 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_1214 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_1229 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1235 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_1256 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1283 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1295 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_1307 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_682 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_688 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_702 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_708 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_726 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_734 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_752 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_758 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_764 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_770 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_849 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_855 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_876 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_882 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_885 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_892 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_902 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_928 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_932 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_935 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_971 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_995 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_1002 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_1013 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_1022 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_1046 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_1052 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_1069 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_1100 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_1106 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_1114 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_1125 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_1129 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_1150 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_1161 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_1167 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_1186 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_1190 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_1198 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_1209 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_1218 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_1224 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_1237 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_1243 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1263 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1275 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_708 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_724 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_730 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_736 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_742 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_779 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_827 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_877 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_883 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_886 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_913 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_917 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_922 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_934 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_941 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_949 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_952 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_971 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_986 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_996 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_1004 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_1012 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_1018 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_1027 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_1034 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_1044 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_1068 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_1074 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_1097 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_1125 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_1131 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_1135 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_1171 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_1181 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_1202 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_1227 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_1251 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_685 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_697 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_710 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_751 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_807 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_825 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_859 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_867 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_902 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_919 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_948 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_976 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_1000 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_1031 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_1055 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_1069 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_1075 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1083 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_1104 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_1112 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_1125 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_1131 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_1137 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_1143 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_1155 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_1161 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_1167 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_1173 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_1181 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_1189 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_1195 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_1201 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_1207 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_1213 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1219 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1231 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1237 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1273 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_713 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_749 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_752 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_762 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_774 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_780 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_786 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_792 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_838 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_848 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_856 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_877 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_902 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_934 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_940 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_946 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_949 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_960 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_979 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_993 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_1030 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_1050 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_1074 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_1080 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_1086 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_1105 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_1114 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_1118 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_1139 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_1145 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_1157 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_1163 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_1191 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_1203 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1209 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1221 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1245 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_758 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_764 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_770 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_792 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_804 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_816 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_824 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_839 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_866 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_870 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_883 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_930 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_934 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_937 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_943 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_968 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_972 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_979 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_990 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_1017 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_1023 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1027 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_1048 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_1069 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_1098 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_1110 ();
 sky130_fd_sc_hd__decap_3 FILLER_181_1117 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_1131 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1145 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_1166 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_1172 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_1187 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_1197 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1209 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_1221 ();
 sky130_fd_sc_hd__decap_3 FILLER_181_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_771 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_777 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_792 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_821 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_849 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_857 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_891 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_903 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_932 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_936 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_940 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_951 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_959 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_966 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_988 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_996 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_1002 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_1014 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_1027 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_1037 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_1041 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_1068 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_1078 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_1086 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_1102 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_1109 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_1117 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_1122 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_1134 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_1159 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_1177 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_1198 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1209 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1221 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1245 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_773 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_779 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_797 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_850 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_856 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_878 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_884 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_907 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_922 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_960 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_967 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_975 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_984 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_991 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_997 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_1023 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_1044 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_1055 ();
 sky130_fd_sc_hd__decap_3 FILLER_183_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_1074 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_1080 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_1088 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_1092 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_1103 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_1128 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_1136 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_1145 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_1157 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_1168 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_1174 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_1186 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_1210 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1216 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_1228 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_779 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_822 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_828 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_835 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_843 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_857 ();
 sky130_fd_sc_hd__decap_3 FILLER_184_865 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_876 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_882 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_903 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_934 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_938 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_942 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_954 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_962 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_968 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_972 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_988 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_994 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1002 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_1008 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_1032 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_1041 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1053 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_1074 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_1081 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_1104 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_1117 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_1131 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_1140 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_1159 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_1165 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1169 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_1178 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_1202 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_1212 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_1221 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1227 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1239 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_1251 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_783 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_822 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_835 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_838 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_854 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_865 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_882 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_895 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_912 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_963 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_969 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_975 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_984 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_995 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_1019 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_1025 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_1052 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_1058 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_1087 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_1098 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_1111 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_1118 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_1121 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_1145 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_1158 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_1168 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_1177 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_1184 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_1190 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_1212 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1218 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_737 ();
 sky130_fd_sc_hd__decap_3 FILLER_186_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_778 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_786 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_792 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_795 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_830 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_840 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_849 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_853 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_862 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_880 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_884 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_895 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_898 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_908 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_912 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_915 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_931 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_939 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_943 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_952 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_970 ();
 sky130_fd_sc_hd__decap_3 FILLER_186_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_990 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_996 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_1005 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_1016 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_1027 ();
 sky130_fd_sc_hd__decap_3 FILLER_186_1033 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_1072 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_1088 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_1103 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_1109 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_1154 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_1166 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_1175 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_1184 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_1192 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_1203 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_1212 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1220 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1232 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1244 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_1256 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_741 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_762 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_792 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_799 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_808 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_848 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_854 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_860 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_867 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_890 ();
 sky130_fd_sc_hd__decap_3 FILLER_187_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_902 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_913 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_920 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_928 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_944 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_950 ();
 sky130_fd_sc_hd__decap_3 FILLER_187_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_975 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_1020 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_1026 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_1036 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_1042 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_1048 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_1062 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_1073 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_1086 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1094 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_1100 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_1111 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_1126 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_1151 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1175 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_1187 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_1197 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_1207 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_777 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_799 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_811 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_836 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_890 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_947 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_964 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_974 ();
 sky130_fd_sc_hd__decap_3 FILLER_188_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_999 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_1005 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_1060 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_1084 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_1090 ();
 sky130_fd_sc_hd__decap_3 FILLER_188_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_1102 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_1128 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_1142 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_1146 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_1153 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_1158 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_1165 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_1190 ();
 sky130_fd_sc_hd__decap_3 FILLER_188_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_797 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_822 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_828 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_839 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_859 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_867 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_919 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_936 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_940 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_943 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_964 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_974 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_1006 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_1018 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_1026 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_1029 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_1053 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_1073 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_1083 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_1106 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_1128 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_1141 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_1168 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_1174 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_1177 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_1189 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_1195 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1217 ();
 sky130_fd_sc_hd__decap_3 FILLER_189_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_772 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_781 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_801 ();
 sky130_fd_sc_hd__decap_3 FILLER_190_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_835 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_842 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_846 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_876 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_883 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_889 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_923 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_940 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_965 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_988 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_994 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_1000 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1008 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_1022 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_1028 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_1045 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_1063 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_1071 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_1075 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_1084 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_1090 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_1107 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_1118 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_1127 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_1133 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_1154 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_1166 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_1176 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_1186 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1192 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_727 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_756 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_768 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_790 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_802 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_814 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_826 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_851 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_864 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_892 ();
 sky130_fd_sc_hd__decap_3 FILLER_191_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_902 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_926 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_950 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_960 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_966 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_977 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_1029 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_1035 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_1042 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_1055 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_1087 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_1100 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_1112 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_1126 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_1134 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_1143 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_1175 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1181 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1193 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1217 ();
 sky130_fd_sc_hd__decap_3 FILLER_191_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_767 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_795 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_810 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_819 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_833 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_854 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_874 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_880 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_886 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_892 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_895 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_929 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_954 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_986 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_992 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1004 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1016 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_1028 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_1041 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_1054 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_1061 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_1067 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_1073 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_1079 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_1086 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_1115 ();
 sky130_fd_sc_hd__decap_3 FILLER_192_1123 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_1154 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_1160 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_1168 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1186 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_1198 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_741 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_759 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_765 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_776 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_814 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_826 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_830 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_848 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_856 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_913 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_922 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_928 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_934 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_940 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_947 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_950 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_973 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1033 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_1045 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_1049 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_1055 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1069 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1081 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_1097 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1106 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_1118 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1121 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1144 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1156 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_1168 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_755 ();
 sky130_fd_sc_hd__decap_3 FILLER_194_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_763 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_771 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_778 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_790 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_822 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_923 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_931 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_934 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_946 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_958 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_873 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_885 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_889 ();
 sky130_fd_sc_hd__decap_8 FILLER_210_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_903 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_907 ();
 sky130_fd_sc_hd__decap_8 FILLER_210_913 ();
 sky130_fd_sc_hd__decap_3 FILLER_210_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_210_937 ();
 sky130_fd_sc_hd__decap_8 FILLER_210_947 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_958 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_964 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_976 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_211_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_26 ();
 sky130_fd_sc_hd__decap_8 FILLER_211_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_73 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_211_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_211_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_211_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_294 ();
 sky130_fd_sc_hd__decap_8 FILLER_211_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_211_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_332 ();
 sky130_fd_sc_hd__decap_8 FILLER_211_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_211_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_211_412 ();
 sky130_fd_sc_hd__decap_8 FILLER_211_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_211_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_538 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_594 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_600 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_604 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_629 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_638 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_651 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_685 ();
 sky130_fd_sc_hd__decap_8 FILLER_211_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_706 ();
 sky130_fd_sc_hd__decap_8 FILLER_211_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_726 ();
 sky130_fd_sc_hd__decap_8 FILLER_211_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_762 ();
 sky130_fd_sc_hd__decap_8 FILLER_211_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_782 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_791 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_803 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_808 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_211_846 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_854 ();
 sky130_fd_sc_hd__decap_8 FILLER_211_860 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_877 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_894 ();
 sky130_fd_sc_hd__decap_8 FILLER_211_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_905 ();
 sky130_fd_sc_hd__decap_8 FILLER_211_911 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_211_931 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_939 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_951 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_957 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_962 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_991 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_995 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1014 ();
 sky130_fd_sc_hd__decap_8 FILLER_211_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_1034 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1046 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_1058 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1071 ();
 sky130_fd_sc_hd__decap_8 FILLER_211_1083 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1098 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_1110 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_1114 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_1145 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_211_1154 ();
 sky130_fd_sc_hd__decap_8 FILLER_211_1165 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1177 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_1189 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_1195 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_1203 ();
 sky130_fd_sc_hd__decap_8 FILLER_211_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1216 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_1228 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1233 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_1245 ();
 sky130_fd_sc_hd__decap_8 FILLER_211_1250 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_1258 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1267 ();
 sky130_fd_sc_hd__decap_8 FILLER_211_1279 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_1287 ();
 sky130_fd_sc_hd__decap_8 FILLER_211_1289 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_1297 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1301 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_1313 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1322 ();
 sky130_fd_sc_hd__decap_8 FILLER_211_1334 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_1342 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1352 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_1364 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1385 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_1397 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_1401 ();
 sky130_fd_sc_hd__decap_8 FILLER_211_1406 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_1414 ();
 sky130_fd_sc_hd__decap_8 FILLER_211_1420 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1429 ();
 sky130_fd_sc_hd__decap_8 FILLER_211_1441 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_1449 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_1454 ();
 sky130_fd_sc_hd__decap_8 FILLER_211_1457 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_1465 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1471 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1485 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_1497 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_1501 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_1511 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1522 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_1534 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1556 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1574 ();
 sky130_fd_sc_hd__decap_8 FILLER_211_1586 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_1594 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_1597 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_1603 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1607 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_1619 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_1623 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1630 ();
 sky130_fd_sc_hd__decap_8 FILLER_211_1642 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_1650 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1658 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_1670 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_1675 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1693 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_1705 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_1709 ();
 sky130_fd_sc_hd__decap_8 FILLER_211_1714 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_1722 ();
 sky130_fd_sc_hd__decap_8 FILLER_211_1726 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_1734 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1737 ();
 sky130_fd_sc_hd__decap_8 FILLER_211_1749 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_1760 ();
 sky130_fd_sc_hd__decap_8 FILLER_211_1765 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_1773 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1777 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1793 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_1805 ();
 sky130_fd_sc_hd__decap_8 FILLER_211_1811 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_1819 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1828 ();
 sky130_fd_sc_hd__decap_8 FILLER_211_1840 ();
 sky130_fd_sc_hd__decap_8 FILLER_211_1849 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_1857 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1862 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_1874 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1882 ();
 sky130_fd_sc_hd__decap_8 FILLER_211_1894 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_1902 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_1905 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_1909 ();
 sky130_fd_sc_hd__decap_8 FILLER_211_1913 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_1921 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_1927 ();
 assign io_oeb[0] = net264;
 assign io_oeb[10] = net274;
 assign io_oeb[11] = net275;
 assign io_oeb[12] = net276;
 assign io_oeb[13] = net277;
 assign io_oeb[14] = net278;
 assign io_oeb[15] = net279;
 assign io_oeb[16] = net63;
 assign io_oeb[19] = net280;
 assign io_oeb[1] = net265;
 assign io_oeb[20] = net64;
 assign io_oeb[21] = net281;
 assign io_oeb[22] = net282;
 assign io_oeb[23] = net283;
 assign io_oeb[24] = net284;
 assign io_oeb[25] = net285;
 assign io_oeb[26] = net286;
 assign io_oeb[27] = net287;
 assign io_oeb[28] = net288;
 assign io_oeb[29] = net289;
 assign io_oeb[2] = net266;
 assign io_oeb[30] = net290;
 assign io_oeb[31] = net291;
 assign io_oeb[32] = net292;
 assign io_oeb[33] = net293;
 assign io_oeb[34] = net294;
 assign io_oeb[35] = net295;
 assign io_oeb[36] = net296;
 assign io_oeb[37] = net297;
 assign io_oeb[3] = net267;
 assign io_oeb[4] = net268;
 assign io_oeb[5] = net269;
 assign io_oeb[6] = net270;
 assign io_oeb[7] = net271;
 assign io_oeb[8] = net272;
 assign io_oeb[9] = net273;
 assign io_out[0] = net65;
 assign io_out[10] = net75;
 assign io_out[11] = net76;
 assign io_out[12] = net77;
 assign io_out[13] = net78;
 assign io_out[14] = net79;
 assign io_out[15] = net80;
 assign io_out[19] = net81;
 assign io_out[1] = net66;
 assign io_out[21] = net82;
 assign io_out[22] = net83;
 assign io_out[23] = net84;
 assign io_out[24] = net85;
 assign io_out[25] = net86;
 assign io_out[26] = net87;
 assign io_out[27] = net88;
 assign io_out[28] = net89;
 assign io_out[29] = net90;
 assign io_out[2] = net67;
 assign io_out[30] = net91;
 assign io_out[31] = net92;
 assign io_out[32] = net93;
 assign io_out[33] = net94;
 assign io_out[34] = net95;
 assign io_out[35] = net96;
 assign io_out[36] = net97;
 assign io_out[37] = net98;
 assign io_out[3] = net68;
 assign io_out[4] = net69;
 assign io_out[5] = net70;
 assign io_out[6] = net71;
 assign io_out[7] = net72;
 assign io_out[8] = net73;
 assign io_out[9] = net74;
 assign irq[0] = net99;
 assign irq[1] = net100;
 assign irq[2] = net101;
 assign la_data_out[0] = net102;
 assign la_data_out[100] = net202;
 assign la_data_out[101] = net203;
 assign la_data_out[102] = net204;
 assign la_data_out[103] = net205;
 assign la_data_out[104] = net206;
 assign la_data_out[105] = net207;
 assign la_data_out[106] = net208;
 assign la_data_out[107] = net209;
 assign la_data_out[108] = net210;
 assign la_data_out[109] = net211;
 assign la_data_out[10] = net112;
 assign la_data_out[110] = net212;
 assign la_data_out[111] = net213;
 assign la_data_out[112] = net214;
 assign la_data_out[113] = net215;
 assign la_data_out[114] = net216;
 assign la_data_out[115] = net217;
 assign la_data_out[116] = net218;
 assign la_data_out[117] = net219;
 assign la_data_out[118] = net220;
 assign la_data_out[119] = net221;
 assign la_data_out[11] = net113;
 assign la_data_out[120] = net222;
 assign la_data_out[121] = net223;
 assign la_data_out[122] = net224;
 assign la_data_out[123] = net225;
 assign la_data_out[124] = net226;
 assign la_data_out[125] = net227;
 assign la_data_out[126] = net228;
 assign la_data_out[127] = net229;
 assign la_data_out[12] = net114;
 assign la_data_out[13] = net115;
 assign la_data_out[14] = net116;
 assign la_data_out[15] = net117;
 assign la_data_out[16] = net118;
 assign la_data_out[17] = net119;
 assign la_data_out[18] = net120;
 assign la_data_out[19] = net121;
 assign la_data_out[1] = net103;
 assign la_data_out[20] = net122;
 assign la_data_out[21] = net123;
 assign la_data_out[22] = net124;
 assign la_data_out[23] = net125;
 assign la_data_out[24] = net126;
 assign la_data_out[25] = net127;
 assign la_data_out[26] = net128;
 assign la_data_out[27] = net129;
 assign la_data_out[28] = net130;
 assign la_data_out[29] = net131;
 assign la_data_out[2] = net104;
 assign la_data_out[30] = net132;
 assign la_data_out[31] = net133;
 assign la_data_out[32] = net134;
 assign la_data_out[33] = net135;
 assign la_data_out[34] = net136;
 assign la_data_out[35] = net137;
 assign la_data_out[36] = net138;
 assign la_data_out[37] = net139;
 assign la_data_out[38] = net140;
 assign la_data_out[39] = net141;
 assign la_data_out[3] = net105;
 assign la_data_out[40] = net142;
 assign la_data_out[41] = net143;
 assign la_data_out[42] = net144;
 assign la_data_out[43] = net145;
 assign la_data_out[44] = net146;
 assign la_data_out[45] = net147;
 assign la_data_out[46] = net148;
 assign la_data_out[47] = net149;
 assign la_data_out[48] = net150;
 assign la_data_out[49] = net151;
 assign la_data_out[4] = net106;
 assign la_data_out[50] = net152;
 assign la_data_out[51] = net153;
 assign la_data_out[52] = net154;
 assign la_data_out[53] = net155;
 assign la_data_out[54] = net156;
 assign la_data_out[55] = net157;
 assign la_data_out[56] = net158;
 assign la_data_out[57] = net159;
 assign la_data_out[58] = net160;
 assign la_data_out[59] = net161;
 assign la_data_out[5] = net107;
 assign la_data_out[60] = net162;
 assign la_data_out[61] = net163;
 assign la_data_out[62] = net164;
 assign la_data_out[63] = net165;
 assign la_data_out[64] = net166;
 assign la_data_out[65] = net167;
 assign la_data_out[66] = net168;
 assign la_data_out[67] = net169;
 assign la_data_out[68] = net170;
 assign la_data_out[69] = net171;
 assign la_data_out[6] = net108;
 assign la_data_out[70] = net172;
 assign la_data_out[71] = net173;
 assign la_data_out[72] = net174;
 assign la_data_out[73] = net175;
 assign la_data_out[74] = net176;
 assign la_data_out[75] = net177;
 assign la_data_out[76] = net178;
 assign la_data_out[77] = net179;
 assign la_data_out[78] = net180;
 assign la_data_out[79] = net181;
 assign la_data_out[7] = net109;
 assign la_data_out[80] = net182;
 assign la_data_out[81] = net183;
 assign la_data_out[82] = net184;
 assign la_data_out[83] = net185;
 assign la_data_out[84] = net186;
 assign la_data_out[85] = net187;
 assign la_data_out[86] = net188;
 assign la_data_out[87] = net189;
 assign la_data_out[88] = net190;
 assign la_data_out[89] = net191;
 assign la_data_out[8] = net110;
 assign la_data_out[90] = net192;
 assign la_data_out[91] = net193;
 assign la_data_out[92] = net194;
 assign la_data_out[93] = net195;
 assign la_data_out[94] = net196;
 assign la_data_out[95] = net197;
 assign la_data_out[96] = net198;
 assign la_data_out[97] = net199;
 assign la_data_out[98] = net200;
 assign la_data_out[99] = net201;
 assign la_data_out[9] = net111;
 assign wbs_ack_o = net230;
 assign wbs_dat_o[0] = net231;
 assign wbs_dat_o[10] = net241;
 assign wbs_dat_o[11] = net242;
 assign wbs_dat_o[12] = net243;
 assign wbs_dat_o[13] = net244;
 assign wbs_dat_o[14] = net245;
 assign wbs_dat_o[15] = net246;
 assign wbs_dat_o[16] = net247;
 assign wbs_dat_o[17] = net248;
 assign wbs_dat_o[18] = net249;
 assign wbs_dat_o[19] = net250;
 assign wbs_dat_o[1] = net232;
 assign wbs_dat_o[20] = net251;
 assign wbs_dat_o[21] = net252;
 assign wbs_dat_o[22] = net253;
 assign wbs_dat_o[23] = net254;
 assign wbs_dat_o[24] = net255;
 assign wbs_dat_o[25] = net256;
 assign wbs_dat_o[26] = net257;
 assign wbs_dat_o[27] = net258;
 assign wbs_dat_o[28] = net259;
 assign wbs_dat_o[29] = net260;
 assign wbs_dat_o[2] = net233;
 assign wbs_dat_o[30] = net261;
 assign wbs_dat_o[31] = net262;
 assign wbs_dat_o[3] = net234;
 assign wbs_dat_o[4] = net235;
 assign wbs_dat_o[5] = net236;
 assign wbs_dat_o[6] = net237;
 assign wbs_dat_o[7] = net238;
 assign wbs_dat_o[8] = net239;
 assign wbs_dat_o[9] = net240;
endmodule

